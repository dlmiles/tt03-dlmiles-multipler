
`define	IMPL_TWOS		1
