// headline config
`define X_WIDTH		7
`define Y_WIDTH		7
`define P_WIDTH		14
`define	S_WIDTH		0

// wire [7:0] io_in, interface
`define I_CLK_BITID	0
`define I0_X_BITID	1
`define I1_Y_BITID	1

// wire [7:0] io_out, interface
`define O0_P_LSB_BITID	1
`define O1_P_MSB_BITID	1
