
`define	IMPL_MULU_M3Q3		1
