
`define	IMPL_HALFADDER		1
