// headline config
`define WIDTH		1

// wire [7:0] io_in, interface
`define I_CLK_BITID	0
`define I_RST_BITID	1
`define I_A_BITID	2
`define I_B_BITID	3
`define I_Y_BITID	4

// wire [7:0] io_out, interface
`define O_CARRY_BITID	6
`define O_SUM_BITID	7
