
`define	IMPL_ONES		1
