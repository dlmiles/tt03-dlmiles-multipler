
`define	IMPL_NEGEDGE_CARRY_LOOK_AHEAD		1
