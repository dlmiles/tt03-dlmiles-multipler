// headline config
`define WIDTH		7

// wire [7:0] io_in, interface
`define I_CLK_BITID	0
`define I0_A_BITID	1
`define I0_B_BITID	1

// wire [7:0] io_out, interface
`define O_CARRY_BITID	0
`define O_SUM_BITID	1
