
`define	IMPL_MULU_X2Y2		1
