
`define	IMPL_MULU_M2Q2		1
