`default_nettype none
`timescale 1ns/1ps

/*
this testbench just instantiates the module and makes some convenient wires
that can be driven / tested by the cocotb test.py
*/

module tb_muls_x3y3 (
    // testbench is controlled by test.py
    input clk,
    input rst,
    input [2:0] x,
    input [2:0] y,
    output [5:0] p,
    output s,
    output rdy
);

    // this part dumps the trace to a vcd file that can be viewed with GTKWave
    initial begin
        $dumpfile ("tb_muls_x3y3.vcd");
        $dumpvars (0, tb_muls_x3y3);
        #1;
    end

    // wire up the inputs and outputs
    wire [7:0] inputs = {{y}, {x}, rst, clk};
    wire [7:0] outputs;
    assign p = outputs[5:0];
    assign s = outputs[6];
    assign rdy = outputs[7];

    // instantiate the DUT
    muls_x3y3 multipler_signed_x3y3(
`ifdef GL_TEST
        .vccd1( 1'b1),
        .vssd1( 1'b0),
`endif
        .io_in  (inputs),
        .io_out (outputs)
    );

endmodule
