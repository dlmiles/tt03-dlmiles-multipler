
`define	IMPL_MULS_X3Y3		1
