// headline config
`define X_WIDTH		3
`define Y_WIDTH		3
`define P_WIDTH		6
`define S_WIDTH		1

// wire [7:0] io_in, interface
`define I_CLK_BITID	0
`define I_RST_BITID	1
`define I_X_BITID	2
`define I_Y_BITID	5

// wire [7:0] io_out, interface
`define O_P_BITID	0
`define O_SIGN_BITID	6
`define O_READY_BITID	7
