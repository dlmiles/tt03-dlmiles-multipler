
`define	IMPL_FULLADDER		1
