
`define	IMPL_CARRY_LOOK_AHEAD		1
