// headline config
`define X_WIDTH		2
`define Y_WIDTH		2
`define P_WIDTH		4
`define	S_WIDTH		0

// wire [7:0] io_in, interface
`define I_CLK_BITID	0
`define I_RST_BITID	1
`define I_X_BITID	2
`define I_Y_BITID	4

// wire [7:0] io_out, interface
`define O_P_BITID	0
`define O_SIGN_BITID	6
`define O_READY_BITID	7
