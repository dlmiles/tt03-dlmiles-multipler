
`define	IMPL_MULU_X3Y3		1
