`default_nettype none

`include "global.vh"
`include "config.vh"    // mulu_m7q7.vh

// Unsigned Multipler, X width 2, Y width 2, making P result width 4
module mulu_m7q7 (
    input	[`X_WIDTH-1:0]	m,
    input	[`Y_WIDTH-1:0]	q,

    output reg	[`P_WIDTH-1:0]	p
`ifdef HAS_SIGN
    , output			s
`endif
`ifdef HAS_READY
    , output			rdy
`endif
);

    localparam X_WIDTH = `X_WIDTH;
    localparam Y_WIDTH = `Y_WIDTH;
    localparam P_WIDTH = `P_WIDTH;

`ifdef HAS_SIGN
    // sign bit
    assign s = m[X_WIDTH-1] ^ q[Y_WIDTH-1];
`endif
`ifdef HAS_READY
    // always ready
    assign rdy = `READY_TRUE;
`endif

    /////// PARTIAL PRODUCTS

    // This method is better for working when X_WIDTH != Y_WIDTH
    wire [Y_WIDTH-1:0] pp [X_WIDTH-1:0];

    genvar ppiq;
    genvar ppim;
    generate //: genpp
        for (ppiq = 0; ppiq < Y_WIDTH; ppiq = ppiq + 1) begin		// loop 7 times, from 0
            // If X_WIDTH == Y_WIDTH then this for loop below means:
            // pp[iq][X_WIDTH-1:0] = m[X_WIDTH-1:0] & {X_WIDTH{q[ppiq]}}
            for(ppim = 0; ppim < X_WIDTH; ppim = ppim + 1) begin	// loop 7 times, from 0
                assign pp[ppiq][ppim] = m[ppim] & q[ppiq];
            end
        end
    endgenerate
    
    wire [`P_WIDTH-1:0] mq = {m,q};

    always_comb begin
        case (mq)
            {7'd0,7'd0}:		p = 14'd0;
            {7'd0,7'd1}:		p = 14'd0;
            {7'd0,7'd2}:		p = 14'd0;
            {7'd0,7'd3}:		p = 14'd0;
            {7'd0,7'd4}:		p = 14'd0;
            {7'd0,7'd5}:		p = 14'd0;
            {7'd0,7'd6}:		p = 14'd0;
            {7'd0,7'd7}:		p = 14'd0;
            {7'd0,7'd8}:		p = 14'd0;
            {7'd0,7'd9}:		p = 14'd0;
            {7'd0,7'd10}:		p = 14'd0;
            {7'd0,7'd11}:		p = 14'd0;
            {7'd0,7'd12}:		p = 14'd0;
            {7'd0,7'd13}:		p = 14'd0;
            {7'd0,7'd14}:		p = 14'd0;
            {7'd0,7'd15}:		p = 14'd0;
            {7'd0,7'd16}:		p = 14'd0;
            {7'd0,7'd17}:		p = 14'd0;
            {7'd0,7'd18}:		p = 14'd0;
            {7'd0,7'd19}:		p = 14'd0;
            {7'd0,7'd20}:		p = 14'd0;
            {7'd0,7'd21}:		p = 14'd0;
            {7'd0,7'd22}:		p = 14'd0;
            {7'd0,7'd23}:		p = 14'd0;
            {7'd0,7'd24}:		p = 14'd0;
            {7'd0,7'd25}:		p = 14'd0;
            {7'd0,7'd26}:		p = 14'd0;
            {7'd0,7'd27}:		p = 14'd0;
            {7'd0,7'd28}:		p = 14'd0;
            {7'd0,7'd29}:		p = 14'd0;
            {7'd0,7'd30}:		p = 14'd0;
            {7'd0,7'd31}:		p = 14'd0;
            {7'd0,7'd32}:		p = 14'd0;
            {7'd0,7'd33}:		p = 14'd0;
            {7'd0,7'd34}:		p = 14'd0;
            {7'd0,7'd35}:		p = 14'd0;
            {7'd0,7'd36}:		p = 14'd0;
            {7'd0,7'd37}:		p = 14'd0;
            {7'd0,7'd38}:		p = 14'd0;
            {7'd0,7'd39}:		p = 14'd0;
            {7'd0,7'd40}:		p = 14'd0;
            {7'd0,7'd41}:		p = 14'd0;
            {7'd0,7'd42}:		p = 14'd0;
            {7'd0,7'd43}:		p = 14'd0;
            {7'd0,7'd44}:		p = 14'd0;
            {7'd0,7'd45}:		p = 14'd0;
            {7'd0,7'd46}:		p = 14'd0;
            {7'd0,7'd47}:		p = 14'd0;
            {7'd0,7'd48}:		p = 14'd0;
            {7'd0,7'd49}:		p = 14'd0;
            {7'd0,7'd50}:		p = 14'd0;
            {7'd0,7'd51}:		p = 14'd0;
            {7'd0,7'd52}:		p = 14'd0;
            {7'd0,7'd53}:		p = 14'd0;
            {7'd0,7'd54}:		p = 14'd0;
            {7'd0,7'd55}:		p = 14'd0;
            {7'd0,7'd56}:		p = 14'd0;
            {7'd0,7'd57}:		p = 14'd0;
            {7'd0,7'd58}:		p = 14'd0;
            {7'd0,7'd59}:		p = 14'd0;
            {7'd0,7'd60}:		p = 14'd0;
            {7'd0,7'd61}:		p = 14'd0;
            {7'd0,7'd62}:		p = 14'd0;
            {7'd0,7'd63}:		p = 14'd0;
            {7'd0,7'd64}:		p = 14'd0;
            {7'd0,7'd65}:		p = 14'd0;
            {7'd0,7'd66}:		p = 14'd0;
            {7'd0,7'd67}:		p = 14'd0;
            {7'd0,7'd68}:		p = 14'd0;
            {7'd0,7'd69}:		p = 14'd0;
            {7'd0,7'd70}:		p = 14'd0;
            {7'd0,7'd71}:		p = 14'd0;
            {7'd0,7'd72}:		p = 14'd0;
            {7'd0,7'd73}:		p = 14'd0;
            {7'd0,7'd74}:		p = 14'd0;
            {7'd0,7'd75}:		p = 14'd0;
            {7'd0,7'd76}:		p = 14'd0;
            {7'd0,7'd77}:		p = 14'd0;
            {7'd0,7'd78}:		p = 14'd0;
            {7'd0,7'd79}:		p = 14'd0;
            {7'd0,7'd80}:		p = 14'd0;
            {7'd0,7'd81}:		p = 14'd0;
            {7'd0,7'd82}:		p = 14'd0;
            {7'd0,7'd83}:		p = 14'd0;
            {7'd0,7'd84}:		p = 14'd0;
            {7'd0,7'd85}:		p = 14'd0;
            {7'd0,7'd86}:		p = 14'd0;
            {7'd0,7'd87}:		p = 14'd0;
            {7'd0,7'd88}:		p = 14'd0;
            {7'd0,7'd89}:		p = 14'd0;
            {7'd0,7'd90}:		p = 14'd0;
            {7'd0,7'd91}:		p = 14'd0;
            {7'd0,7'd92}:		p = 14'd0;
            {7'd0,7'd93}:		p = 14'd0;
            {7'd0,7'd94}:		p = 14'd0;
            {7'd0,7'd95}:		p = 14'd0;
            {7'd0,7'd96}:		p = 14'd0;
            {7'd0,7'd97}:		p = 14'd0;
            {7'd0,7'd98}:		p = 14'd0;
            {7'd0,7'd99}:		p = 14'd0;
            {7'd0,7'd100}:		p = 14'd0;
            {7'd0,7'd101}:		p = 14'd0;
            {7'd0,7'd102}:		p = 14'd0;
            {7'd0,7'd103}:		p = 14'd0;
            {7'd0,7'd104}:		p = 14'd0;
            {7'd0,7'd105}:		p = 14'd0;
            {7'd0,7'd106}:		p = 14'd0;
            {7'd0,7'd107}:		p = 14'd0;
            {7'd0,7'd108}:		p = 14'd0;
            {7'd0,7'd109}:		p = 14'd0;
            {7'd0,7'd110}:		p = 14'd0;
            {7'd0,7'd111}:		p = 14'd0;
            {7'd0,7'd112}:		p = 14'd0;
            {7'd0,7'd113}:		p = 14'd0;
            {7'd0,7'd114}:		p = 14'd0;
            {7'd0,7'd115}:		p = 14'd0;
            {7'd0,7'd116}:		p = 14'd0;
            {7'd0,7'd117}:		p = 14'd0;
            {7'd0,7'd118}:		p = 14'd0;
            {7'd0,7'd119}:		p = 14'd0;
            {7'd0,7'd120}:		p = 14'd0;
            {7'd0,7'd121}:		p = 14'd0;
            {7'd0,7'd122}:		p = 14'd0;
            {7'd0,7'd123}:		p = 14'd0;
            {7'd0,7'd124}:		p = 14'd0;
            {7'd0,7'd125}:		p = 14'd0;
            {7'd0,7'd126}:		p = 14'd0;
            {7'd0,7'd127}:		p = 14'd0;
            {7'd1,7'd0}:		p = 14'd0;
            {7'd1,7'd1}:		p = 14'd1;
            {7'd1,7'd2}:		p = 14'd2;
            {7'd1,7'd3}:		p = 14'd3;
            {7'd1,7'd4}:		p = 14'd4;
            {7'd1,7'd5}:		p = 14'd5;
            {7'd1,7'd6}:		p = 14'd6;
            {7'd1,7'd7}:		p = 14'd7;
            {7'd1,7'd8}:		p = 14'd8;
            {7'd1,7'd9}:		p = 14'd9;
            {7'd1,7'd10}:		p = 14'd10;
            {7'd1,7'd11}:		p = 14'd11;
            {7'd1,7'd12}:		p = 14'd12;
            {7'd1,7'd13}:		p = 14'd13;
            {7'd1,7'd14}:		p = 14'd14;
            {7'd1,7'd15}:		p = 14'd15;
            {7'd1,7'd16}:		p = 14'd16;
            {7'd1,7'd17}:		p = 14'd17;
            {7'd1,7'd18}:		p = 14'd18;
            {7'd1,7'd19}:		p = 14'd19;
            {7'd1,7'd20}:		p = 14'd20;
            {7'd1,7'd21}:		p = 14'd21;
            {7'd1,7'd22}:		p = 14'd22;
            {7'd1,7'd23}:		p = 14'd23;
            {7'd1,7'd24}:		p = 14'd24;
            {7'd1,7'd25}:		p = 14'd25;
            {7'd1,7'd26}:		p = 14'd26;
            {7'd1,7'd27}:		p = 14'd27;
            {7'd1,7'd28}:		p = 14'd28;
            {7'd1,7'd29}:		p = 14'd29;
            {7'd1,7'd30}:		p = 14'd30;
            {7'd1,7'd31}:		p = 14'd31;
            {7'd1,7'd32}:		p = 14'd32;
            {7'd1,7'd33}:		p = 14'd33;
            {7'd1,7'd34}:		p = 14'd34;
            {7'd1,7'd35}:		p = 14'd35;
            {7'd1,7'd36}:		p = 14'd36;
            {7'd1,7'd37}:		p = 14'd37;
            {7'd1,7'd38}:		p = 14'd38;
            {7'd1,7'd39}:		p = 14'd39;
            {7'd1,7'd40}:		p = 14'd40;
            {7'd1,7'd41}:		p = 14'd41;
            {7'd1,7'd42}:		p = 14'd42;
            {7'd1,7'd43}:		p = 14'd43;
            {7'd1,7'd44}:		p = 14'd44;
            {7'd1,7'd45}:		p = 14'd45;
            {7'd1,7'd46}:		p = 14'd46;
            {7'd1,7'd47}:		p = 14'd47;
            {7'd1,7'd48}:		p = 14'd48;
            {7'd1,7'd49}:		p = 14'd49;
            {7'd1,7'd50}:		p = 14'd50;
            {7'd1,7'd51}:		p = 14'd51;
            {7'd1,7'd52}:		p = 14'd52;
            {7'd1,7'd53}:		p = 14'd53;
            {7'd1,7'd54}:		p = 14'd54;
            {7'd1,7'd55}:		p = 14'd55;
            {7'd1,7'd56}:		p = 14'd56;
            {7'd1,7'd57}:		p = 14'd57;
            {7'd1,7'd58}:		p = 14'd58;
            {7'd1,7'd59}:		p = 14'd59;
            {7'd1,7'd60}:		p = 14'd60;
            {7'd1,7'd61}:		p = 14'd61;
            {7'd1,7'd62}:		p = 14'd62;
            {7'd1,7'd63}:		p = 14'd63;
            {7'd1,7'd64}:		p = 14'd64;
            {7'd1,7'd65}:		p = 14'd65;
            {7'd1,7'd66}:		p = 14'd66;
            {7'd1,7'd67}:		p = 14'd67;
            {7'd1,7'd68}:		p = 14'd68;
            {7'd1,7'd69}:		p = 14'd69;
            {7'd1,7'd70}:		p = 14'd70;
            {7'd1,7'd71}:		p = 14'd71;
            {7'd1,7'd72}:		p = 14'd72;
            {7'd1,7'd73}:		p = 14'd73;
            {7'd1,7'd74}:		p = 14'd74;
            {7'd1,7'd75}:		p = 14'd75;
            {7'd1,7'd76}:		p = 14'd76;
            {7'd1,7'd77}:		p = 14'd77;
            {7'd1,7'd78}:		p = 14'd78;
            {7'd1,7'd79}:		p = 14'd79;
            {7'd1,7'd80}:		p = 14'd80;
            {7'd1,7'd81}:		p = 14'd81;
            {7'd1,7'd82}:		p = 14'd82;
            {7'd1,7'd83}:		p = 14'd83;
            {7'd1,7'd84}:		p = 14'd84;
            {7'd1,7'd85}:		p = 14'd85;
            {7'd1,7'd86}:		p = 14'd86;
            {7'd1,7'd87}:		p = 14'd87;
            {7'd1,7'd88}:		p = 14'd88;
            {7'd1,7'd89}:		p = 14'd89;
            {7'd1,7'd90}:		p = 14'd90;
            {7'd1,7'd91}:		p = 14'd91;
            {7'd1,7'd92}:		p = 14'd92;
            {7'd1,7'd93}:		p = 14'd93;
            {7'd1,7'd94}:		p = 14'd94;
            {7'd1,7'd95}:		p = 14'd95;
            {7'd1,7'd96}:		p = 14'd96;
            {7'd1,7'd97}:		p = 14'd97;
            {7'd1,7'd98}:		p = 14'd98;
            {7'd1,7'd99}:		p = 14'd99;
            {7'd1,7'd100}:		p = 14'd100;
            {7'd1,7'd101}:		p = 14'd101;
            {7'd1,7'd102}:		p = 14'd102;
            {7'd1,7'd103}:		p = 14'd103;
            {7'd1,7'd104}:		p = 14'd104;
            {7'd1,7'd105}:		p = 14'd105;
            {7'd1,7'd106}:		p = 14'd106;
            {7'd1,7'd107}:		p = 14'd107;
            {7'd1,7'd108}:		p = 14'd108;
            {7'd1,7'd109}:		p = 14'd109;
            {7'd1,7'd110}:		p = 14'd110;
            {7'd1,7'd111}:		p = 14'd111;
            {7'd1,7'd112}:		p = 14'd112;
            {7'd1,7'd113}:		p = 14'd113;
            {7'd1,7'd114}:		p = 14'd114;
            {7'd1,7'd115}:		p = 14'd115;
            {7'd1,7'd116}:		p = 14'd116;
            {7'd1,7'd117}:		p = 14'd117;
            {7'd1,7'd118}:		p = 14'd118;
            {7'd1,7'd119}:		p = 14'd119;
            {7'd1,7'd120}:		p = 14'd120;
            {7'd1,7'd121}:		p = 14'd121;
            {7'd1,7'd122}:		p = 14'd122;
            {7'd1,7'd123}:		p = 14'd123;
            {7'd1,7'd124}:		p = 14'd124;
            {7'd1,7'd125}:		p = 14'd125;
            {7'd1,7'd126}:		p = 14'd126;
            {7'd1,7'd127}:		p = 14'd127;
            {7'd2,7'd0}:		p = 14'd0;
            {7'd2,7'd1}:		p = 14'd2;
            {7'd2,7'd2}:		p = 14'd4;
            {7'd2,7'd3}:		p = 14'd6;
            {7'd2,7'd4}:		p = 14'd8;
            {7'd2,7'd5}:		p = 14'd10;
            {7'd2,7'd6}:		p = 14'd12;
            {7'd2,7'd7}:		p = 14'd14;
            {7'd2,7'd8}:		p = 14'd16;
            {7'd2,7'd9}:		p = 14'd18;
            {7'd2,7'd10}:		p = 14'd20;
            {7'd2,7'd11}:		p = 14'd22;
            {7'd2,7'd12}:		p = 14'd24;
            {7'd2,7'd13}:		p = 14'd26;
            {7'd2,7'd14}:		p = 14'd28;
            {7'd2,7'd15}:		p = 14'd30;
            {7'd2,7'd16}:		p = 14'd32;
            {7'd2,7'd17}:		p = 14'd34;
            {7'd2,7'd18}:		p = 14'd36;
            {7'd2,7'd19}:		p = 14'd38;
            {7'd2,7'd20}:		p = 14'd40;
            {7'd2,7'd21}:		p = 14'd42;
            {7'd2,7'd22}:		p = 14'd44;
            {7'd2,7'd23}:		p = 14'd46;
            {7'd2,7'd24}:		p = 14'd48;
            {7'd2,7'd25}:		p = 14'd50;
            {7'd2,7'd26}:		p = 14'd52;
            {7'd2,7'd27}:		p = 14'd54;
            {7'd2,7'd28}:		p = 14'd56;
            {7'd2,7'd29}:		p = 14'd58;
            {7'd2,7'd30}:		p = 14'd60;
            {7'd2,7'd31}:		p = 14'd62;
            {7'd2,7'd32}:		p = 14'd64;
            {7'd2,7'd33}:		p = 14'd66;
            {7'd2,7'd34}:		p = 14'd68;
            {7'd2,7'd35}:		p = 14'd70;
            {7'd2,7'd36}:		p = 14'd72;
            {7'd2,7'd37}:		p = 14'd74;
            {7'd2,7'd38}:		p = 14'd76;
            {7'd2,7'd39}:		p = 14'd78;
            {7'd2,7'd40}:		p = 14'd80;
            {7'd2,7'd41}:		p = 14'd82;
            {7'd2,7'd42}:		p = 14'd84;
            {7'd2,7'd43}:		p = 14'd86;
            {7'd2,7'd44}:		p = 14'd88;
            {7'd2,7'd45}:		p = 14'd90;
            {7'd2,7'd46}:		p = 14'd92;
            {7'd2,7'd47}:		p = 14'd94;
            {7'd2,7'd48}:		p = 14'd96;
            {7'd2,7'd49}:		p = 14'd98;
            {7'd2,7'd50}:		p = 14'd100;
            {7'd2,7'd51}:		p = 14'd102;
            {7'd2,7'd52}:		p = 14'd104;
            {7'd2,7'd53}:		p = 14'd106;
            {7'd2,7'd54}:		p = 14'd108;
            {7'd2,7'd55}:		p = 14'd110;
            {7'd2,7'd56}:		p = 14'd112;
            {7'd2,7'd57}:		p = 14'd114;
            {7'd2,7'd58}:		p = 14'd116;
            {7'd2,7'd59}:		p = 14'd118;
            {7'd2,7'd60}:		p = 14'd120;
            {7'd2,7'd61}:		p = 14'd122;
            {7'd2,7'd62}:		p = 14'd124;
            {7'd2,7'd63}:		p = 14'd126;
            {7'd2,7'd64}:		p = 14'd128;
            {7'd2,7'd65}:		p = 14'd130;
            {7'd2,7'd66}:		p = 14'd132;
            {7'd2,7'd67}:		p = 14'd134;
            {7'd2,7'd68}:		p = 14'd136;
            {7'd2,7'd69}:		p = 14'd138;
            {7'd2,7'd70}:		p = 14'd140;
            {7'd2,7'd71}:		p = 14'd142;
            {7'd2,7'd72}:		p = 14'd144;
            {7'd2,7'd73}:		p = 14'd146;
            {7'd2,7'd74}:		p = 14'd148;
            {7'd2,7'd75}:		p = 14'd150;
            {7'd2,7'd76}:		p = 14'd152;
            {7'd2,7'd77}:		p = 14'd154;
            {7'd2,7'd78}:		p = 14'd156;
            {7'd2,7'd79}:		p = 14'd158;
            {7'd2,7'd80}:		p = 14'd160;
            {7'd2,7'd81}:		p = 14'd162;
            {7'd2,7'd82}:		p = 14'd164;
            {7'd2,7'd83}:		p = 14'd166;
            {7'd2,7'd84}:		p = 14'd168;
            {7'd2,7'd85}:		p = 14'd170;
            {7'd2,7'd86}:		p = 14'd172;
            {7'd2,7'd87}:		p = 14'd174;
            {7'd2,7'd88}:		p = 14'd176;
            {7'd2,7'd89}:		p = 14'd178;
            {7'd2,7'd90}:		p = 14'd180;
            {7'd2,7'd91}:		p = 14'd182;
            {7'd2,7'd92}:		p = 14'd184;
            {7'd2,7'd93}:		p = 14'd186;
            {7'd2,7'd94}:		p = 14'd188;
            {7'd2,7'd95}:		p = 14'd190;
            {7'd2,7'd96}:		p = 14'd192;
            {7'd2,7'd97}:		p = 14'd194;
            {7'd2,7'd98}:		p = 14'd196;
            {7'd2,7'd99}:		p = 14'd198;
            {7'd2,7'd100}:		p = 14'd200;
            {7'd2,7'd101}:		p = 14'd202;
            {7'd2,7'd102}:		p = 14'd204;
            {7'd2,7'd103}:		p = 14'd206;
            {7'd2,7'd104}:		p = 14'd208;
            {7'd2,7'd105}:		p = 14'd210;
            {7'd2,7'd106}:		p = 14'd212;
            {7'd2,7'd107}:		p = 14'd214;
            {7'd2,7'd108}:		p = 14'd216;
            {7'd2,7'd109}:		p = 14'd218;
            {7'd2,7'd110}:		p = 14'd220;
            {7'd2,7'd111}:		p = 14'd222;
            {7'd2,7'd112}:		p = 14'd224;
            {7'd2,7'd113}:		p = 14'd226;
            {7'd2,7'd114}:		p = 14'd228;
            {7'd2,7'd115}:		p = 14'd230;
            {7'd2,7'd116}:		p = 14'd232;
            {7'd2,7'd117}:		p = 14'd234;
            {7'd2,7'd118}:		p = 14'd236;
            {7'd2,7'd119}:		p = 14'd238;
            {7'd2,7'd120}:		p = 14'd240;
            {7'd2,7'd121}:		p = 14'd242;
            {7'd2,7'd122}:		p = 14'd244;
            {7'd2,7'd123}:		p = 14'd246;
            {7'd2,7'd124}:		p = 14'd248;
            {7'd2,7'd125}:		p = 14'd250;
            {7'd2,7'd126}:		p = 14'd252;
            {7'd2,7'd127}:		p = 14'd254;
            {7'd3,7'd0}:		p = 14'd0;
            {7'd3,7'd1}:		p = 14'd3;
            {7'd3,7'd2}:		p = 14'd6;
            {7'd3,7'd3}:		p = 14'd9;
            {7'd3,7'd4}:		p = 14'd12;
            {7'd3,7'd5}:		p = 14'd15;
            {7'd3,7'd6}:		p = 14'd18;
            {7'd3,7'd7}:		p = 14'd21;
            {7'd3,7'd8}:		p = 14'd24;
            {7'd3,7'd9}:		p = 14'd27;
            {7'd3,7'd10}:		p = 14'd30;
            {7'd3,7'd11}:		p = 14'd33;
            {7'd3,7'd12}:		p = 14'd36;
            {7'd3,7'd13}:		p = 14'd39;
            {7'd3,7'd14}:		p = 14'd42;
            {7'd3,7'd15}:		p = 14'd45;
            {7'd3,7'd16}:		p = 14'd48;
            {7'd3,7'd17}:		p = 14'd51;
            {7'd3,7'd18}:		p = 14'd54;
            {7'd3,7'd19}:		p = 14'd57;
            {7'd3,7'd20}:		p = 14'd60;
            {7'd3,7'd21}:		p = 14'd63;
            {7'd3,7'd22}:		p = 14'd66;
            {7'd3,7'd23}:		p = 14'd69;
            {7'd3,7'd24}:		p = 14'd72;
            {7'd3,7'd25}:		p = 14'd75;
            {7'd3,7'd26}:		p = 14'd78;
            {7'd3,7'd27}:		p = 14'd81;
            {7'd3,7'd28}:		p = 14'd84;
            {7'd3,7'd29}:		p = 14'd87;
            {7'd3,7'd30}:		p = 14'd90;
            {7'd3,7'd31}:		p = 14'd93;
            {7'd3,7'd32}:		p = 14'd96;
            {7'd3,7'd33}:		p = 14'd99;
            {7'd3,7'd34}:		p = 14'd102;
            {7'd3,7'd35}:		p = 14'd105;
            {7'd3,7'd36}:		p = 14'd108;
            {7'd3,7'd37}:		p = 14'd111;
            {7'd3,7'd38}:		p = 14'd114;
            {7'd3,7'd39}:		p = 14'd117;
            {7'd3,7'd40}:		p = 14'd120;
            {7'd3,7'd41}:		p = 14'd123;
            {7'd3,7'd42}:		p = 14'd126;
            {7'd3,7'd43}:		p = 14'd129;
            {7'd3,7'd44}:		p = 14'd132;
            {7'd3,7'd45}:		p = 14'd135;
            {7'd3,7'd46}:		p = 14'd138;
            {7'd3,7'd47}:		p = 14'd141;
            {7'd3,7'd48}:		p = 14'd144;
            {7'd3,7'd49}:		p = 14'd147;
            {7'd3,7'd50}:		p = 14'd150;
            {7'd3,7'd51}:		p = 14'd153;
            {7'd3,7'd52}:		p = 14'd156;
            {7'd3,7'd53}:		p = 14'd159;
            {7'd3,7'd54}:		p = 14'd162;
            {7'd3,7'd55}:		p = 14'd165;
            {7'd3,7'd56}:		p = 14'd168;
            {7'd3,7'd57}:		p = 14'd171;
            {7'd3,7'd58}:		p = 14'd174;
            {7'd3,7'd59}:		p = 14'd177;
            {7'd3,7'd60}:		p = 14'd180;
            {7'd3,7'd61}:		p = 14'd183;
            {7'd3,7'd62}:		p = 14'd186;
            {7'd3,7'd63}:		p = 14'd189;
            {7'd3,7'd64}:		p = 14'd192;
            {7'd3,7'd65}:		p = 14'd195;
            {7'd3,7'd66}:		p = 14'd198;
            {7'd3,7'd67}:		p = 14'd201;
            {7'd3,7'd68}:		p = 14'd204;
            {7'd3,7'd69}:		p = 14'd207;
            {7'd3,7'd70}:		p = 14'd210;
            {7'd3,7'd71}:		p = 14'd213;
            {7'd3,7'd72}:		p = 14'd216;
            {7'd3,7'd73}:		p = 14'd219;
            {7'd3,7'd74}:		p = 14'd222;
            {7'd3,7'd75}:		p = 14'd225;
            {7'd3,7'd76}:		p = 14'd228;
            {7'd3,7'd77}:		p = 14'd231;
            {7'd3,7'd78}:		p = 14'd234;
            {7'd3,7'd79}:		p = 14'd237;
            {7'd3,7'd80}:		p = 14'd240;
            {7'd3,7'd81}:		p = 14'd243;
            {7'd3,7'd82}:		p = 14'd246;
            {7'd3,7'd83}:		p = 14'd249;
            {7'd3,7'd84}:		p = 14'd252;
            {7'd3,7'd85}:		p = 14'd255;
            {7'd3,7'd86}:		p = 14'd258;
            {7'd3,7'd87}:		p = 14'd261;
            {7'd3,7'd88}:		p = 14'd264;
            {7'd3,7'd89}:		p = 14'd267;
            {7'd3,7'd90}:		p = 14'd270;
            {7'd3,7'd91}:		p = 14'd273;
            {7'd3,7'd92}:		p = 14'd276;
            {7'd3,7'd93}:		p = 14'd279;
            {7'd3,7'd94}:		p = 14'd282;
            {7'd3,7'd95}:		p = 14'd285;
            {7'd3,7'd96}:		p = 14'd288;
            {7'd3,7'd97}:		p = 14'd291;
            {7'd3,7'd98}:		p = 14'd294;
            {7'd3,7'd99}:		p = 14'd297;
            {7'd3,7'd100}:		p = 14'd300;
            {7'd3,7'd101}:		p = 14'd303;
            {7'd3,7'd102}:		p = 14'd306;
            {7'd3,7'd103}:		p = 14'd309;
            {7'd3,7'd104}:		p = 14'd312;
            {7'd3,7'd105}:		p = 14'd315;
            {7'd3,7'd106}:		p = 14'd318;
            {7'd3,7'd107}:		p = 14'd321;
            {7'd3,7'd108}:		p = 14'd324;
            {7'd3,7'd109}:		p = 14'd327;
            {7'd3,7'd110}:		p = 14'd330;
            {7'd3,7'd111}:		p = 14'd333;
            {7'd3,7'd112}:		p = 14'd336;
            {7'd3,7'd113}:		p = 14'd339;
            {7'd3,7'd114}:		p = 14'd342;
            {7'd3,7'd115}:		p = 14'd345;
            {7'd3,7'd116}:		p = 14'd348;
            {7'd3,7'd117}:		p = 14'd351;
            {7'd3,7'd118}:		p = 14'd354;
            {7'd3,7'd119}:		p = 14'd357;
            {7'd3,7'd120}:		p = 14'd360;
            {7'd3,7'd121}:		p = 14'd363;
            {7'd3,7'd122}:		p = 14'd366;
            {7'd3,7'd123}:		p = 14'd369;
            {7'd3,7'd124}:		p = 14'd372;
            {7'd3,7'd125}:		p = 14'd375;
            {7'd3,7'd126}:		p = 14'd378;
            {7'd3,7'd127}:		p = 14'd381;
            {7'd4,7'd0}:		p = 14'd0;
            {7'd4,7'd1}:		p = 14'd4;
            {7'd4,7'd2}:		p = 14'd8;
            {7'd4,7'd3}:		p = 14'd12;
            {7'd4,7'd4}:		p = 14'd16;
            {7'd4,7'd5}:		p = 14'd20;
            {7'd4,7'd6}:		p = 14'd24;
            {7'd4,7'd7}:		p = 14'd28;
            {7'd4,7'd8}:		p = 14'd32;
            {7'd4,7'd9}:		p = 14'd36;
            {7'd4,7'd10}:		p = 14'd40;
            {7'd4,7'd11}:		p = 14'd44;
            {7'd4,7'd12}:		p = 14'd48;
            {7'd4,7'd13}:		p = 14'd52;
            {7'd4,7'd14}:		p = 14'd56;
            {7'd4,7'd15}:		p = 14'd60;
            {7'd4,7'd16}:		p = 14'd64;
            {7'd4,7'd17}:		p = 14'd68;
            {7'd4,7'd18}:		p = 14'd72;
            {7'd4,7'd19}:		p = 14'd76;
            {7'd4,7'd20}:		p = 14'd80;
            {7'd4,7'd21}:		p = 14'd84;
            {7'd4,7'd22}:		p = 14'd88;
            {7'd4,7'd23}:		p = 14'd92;
            {7'd4,7'd24}:		p = 14'd96;
            {7'd4,7'd25}:		p = 14'd100;
            {7'd4,7'd26}:		p = 14'd104;
            {7'd4,7'd27}:		p = 14'd108;
            {7'd4,7'd28}:		p = 14'd112;
            {7'd4,7'd29}:		p = 14'd116;
            {7'd4,7'd30}:		p = 14'd120;
            {7'd4,7'd31}:		p = 14'd124;
            {7'd4,7'd32}:		p = 14'd128;
            {7'd4,7'd33}:		p = 14'd132;
            {7'd4,7'd34}:		p = 14'd136;
            {7'd4,7'd35}:		p = 14'd140;
            {7'd4,7'd36}:		p = 14'd144;
            {7'd4,7'd37}:		p = 14'd148;
            {7'd4,7'd38}:		p = 14'd152;
            {7'd4,7'd39}:		p = 14'd156;
            {7'd4,7'd40}:		p = 14'd160;
            {7'd4,7'd41}:		p = 14'd164;
            {7'd4,7'd42}:		p = 14'd168;
            {7'd4,7'd43}:		p = 14'd172;
            {7'd4,7'd44}:		p = 14'd176;
            {7'd4,7'd45}:		p = 14'd180;
            {7'd4,7'd46}:		p = 14'd184;
            {7'd4,7'd47}:		p = 14'd188;
            {7'd4,7'd48}:		p = 14'd192;
            {7'd4,7'd49}:		p = 14'd196;
            {7'd4,7'd50}:		p = 14'd200;
            {7'd4,7'd51}:		p = 14'd204;
            {7'd4,7'd52}:		p = 14'd208;
            {7'd4,7'd53}:		p = 14'd212;
            {7'd4,7'd54}:		p = 14'd216;
            {7'd4,7'd55}:		p = 14'd220;
            {7'd4,7'd56}:		p = 14'd224;
            {7'd4,7'd57}:		p = 14'd228;
            {7'd4,7'd58}:		p = 14'd232;
            {7'd4,7'd59}:		p = 14'd236;
            {7'd4,7'd60}:		p = 14'd240;
            {7'd4,7'd61}:		p = 14'd244;
            {7'd4,7'd62}:		p = 14'd248;
            {7'd4,7'd63}:		p = 14'd252;
            {7'd4,7'd64}:		p = 14'd256;
            {7'd4,7'd65}:		p = 14'd260;
            {7'd4,7'd66}:		p = 14'd264;
            {7'd4,7'd67}:		p = 14'd268;
            {7'd4,7'd68}:		p = 14'd272;
            {7'd4,7'd69}:		p = 14'd276;
            {7'd4,7'd70}:		p = 14'd280;
            {7'd4,7'd71}:		p = 14'd284;
            {7'd4,7'd72}:		p = 14'd288;
            {7'd4,7'd73}:		p = 14'd292;
            {7'd4,7'd74}:		p = 14'd296;
            {7'd4,7'd75}:		p = 14'd300;
            {7'd4,7'd76}:		p = 14'd304;
            {7'd4,7'd77}:		p = 14'd308;
            {7'd4,7'd78}:		p = 14'd312;
            {7'd4,7'd79}:		p = 14'd316;
            {7'd4,7'd80}:		p = 14'd320;
            {7'd4,7'd81}:		p = 14'd324;
            {7'd4,7'd82}:		p = 14'd328;
            {7'd4,7'd83}:		p = 14'd332;
            {7'd4,7'd84}:		p = 14'd336;
            {7'd4,7'd85}:		p = 14'd340;
            {7'd4,7'd86}:		p = 14'd344;
            {7'd4,7'd87}:		p = 14'd348;
            {7'd4,7'd88}:		p = 14'd352;
            {7'd4,7'd89}:		p = 14'd356;
            {7'd4,7'd90}:		p = 14'd360;
            {7'd4,7'd91}:		p = 14'd364;
            {7'd4,7'd92}:		p = 14'd368;
            {7'd4,7'd93}:		p = 14'd372;
            {7'd4,7'd94}:		p = 14'd376;
            {7'd4,7'd95}:		p = 14'd380;
            {7'd4,7'd96}:		p = 14'd384;
            {7'd4,7'd97}:		p = 14'd388;
            {7'd4,7'd98}:		p = 14'd392;
            {7'd4,7'd99}:		p = 14'd396;
            {7'd4,7'd100}:		p = 14'd400;
            {7'd4,7'd101}:		p = 14'd404;
            {7'd4,7'd102}:		p = 14'd408;
            {7'd4,7'd103}:		p = 14'd412;
            {7'd4,7'd104}:		p = 14'd416;
            {7'd4,7'd105}:		p = 14'd420;
            {7'd4,7'd106}:		p = 14'd424;
            {7'd4,7'd107}:		p = 14'd428;
            {7'd4,7'd108}:		p = 14'd432;
            {7'd4,7'd109}:		p = 14'd436;
            {7'd4,7'd110}:		p = 14'd440;
            {7'd4,7'd111}:		p = 14'd444;
            {7'd4,7'd112}:		p = 14'd448;
            {7'd4,7'd113}:		p = 14'd452;
            {7'd4,7'd114}:		p = 14'd456;
            {7'd4,7'd115}:		p = 14'd460;
            {7'd4,7'd116}:		p = 14'd464;
            {7'd4,7'd117}:		p = 14'd468;
            {7'd4,7'd118}:		p = 14'd472;
            {7'd4,7'd119}:		p = 14'd476;
            {7'd4,7'd120}:		p = 14'd480;
            {7'd4,7'd121}:		p = 14'd484;
            {7'd4,7'd122}:		p = 14'd488;
            {7'd4,7'd123}:		p = 14'd492;
            {7'd4,7'd124}:		p = 14'd496;
            {7'd4,7'd125}:		p = 14'd500;
            {7'd4,7'd126}:		p = 14'd504;
            {7'd4,7'd127}:		p = 14'd508;
            {7'd5,7'd0}:		p = 14'd0;
            {7'd5,7'd1}:		p = 14'd5;
            {7'd5,7'd2}:		p = 14'd10;
            {7'd5,7'd3}:		p = 14'd15;
            {7'd5,7'd4}:		p = 14'd20;
            {7'd5,7'd5}:		p = 14'd25;
            {7'd5,7'd6}:		p = 14'd30;
            {7'd5,7'd7}:		p = 14'd35;
            {7'd5,7'd8}:		p = 14'd40;
            {7'd5,7'd9}:		p = 14'd45;
            {7'd5,7'd10}:		p = 14'd50;
            {7'd5,7'd11}:		p = 14'd55;
            {7'd5,7'd12}:		p = 14'd60;
            {7'd5,7'd13}:		p = 14'd65;
            {7'd5,7'd14}:		p = 14'd70;
            {7'd5,7'd15}:		p = 14'd75;
            {7'd5,7'd16}:		p = 14'd80;
            {7'd5,7'd17}:		p = 14'd85;
            {7'd5,7'd18}:		p = 14'd90;
            {7'd5,7'd19}:		p = 14'd95;
            {7'd5,7'd20}:		p = 14'd100;
            {7'd5,7'd21}:		p = 14'd105;
            {7'd5,7'd22}:		p = 14'd110;
            {7'd5,7'd23}:		p = 14'd115;
            {7'd5,7'd24}:		p = 14'd120;
            {7'd5,7'd25}:		p = 14'd125;
            {7'd5,7'd26}:		p = 14'd130;
            {7'd5,7'd27}:		p = 14'd135;
            {7'd5,7'd28}:		p = 14'd140;
            {7'd5,7'd29}:		p = 14'd145;
            {7'd5,7'd30}:		p = 14'd150;
            {7'd5,7'd31}:		p = 14'd155;
            {7'd5,7'd32}:		p = 14'd160;
            {7'd5,7'd33}:		p = 14'd165;
            {7'd5,7'd34}:		p = 14'd170;
            {7'd5,7'd35}:		p = 14'd175;
            {7'd5,7'd36}:		p = 14'd180;
            {7'd5,7'd37}:		p = 14'd185;
            {7'd5,7'd38}:		p = 14'd190;
            {7'd5,7'd39}:		p = 14'd195;
            {7'd5,7'd40}:		p = 14'd200;
            {7'd5,7'd41}:		p = 14'd205;
            {7'd5,7'd42}:		p = 14'd210;
            {7'd5,7'd43}:		p = 14'd215;
            {7'd5,7'd44}:		p = 14'd220;
            {7'd5,7'd45}:		p = 14'd225;
            {7'd5,7'd46}:		p = 14'd230;
            {7'd5,7'd47}:		p = 14'd235;
            {7'd5,7'd48}:		p = 14'd240;
            {7'd5,7'd49}:		p = 14'd245;
            {7'd5,7'd50}:		p = 14'd250;
            {7'd5,7'd51}:		p = 14'd255;
            {7'd5,7'd52}:		p = 14'd260;
            {7'd5,7'd53}:		p = 14'd265;
            {7'd5,7'd54}:		p = 14'd270;
            {7'd5,7'd55}:		p = 14'd275;
            {7'd5,7'd56}:		p = 14'd280;
            {7'd5,7'd57}:		p = 14'd285;
            {7'd5,7'd58}:		p = 14'd290;
            {7'd5,7'd59}:		p = 14'd295;
            {7'd5,7'd60}:		p = 14'd300;
            {7'd5,7'd61}:		p = 14'd305;
            {7'd5,7'd62}:		p = 14'd310;
            {7'd5,7'd63}:		p = 14'd315;
            {7'd5,7'd64}:		p = 14'd320;
            {7'd5,7'd65}:		p = 14'd325;
            {7'd5,7'd66}:		p = 14'd330;
            {7'd5,7'd67}:		p = 14'd335;
            {7'd5,7'd68}:		p = 14'd340;
            {7'd5,7'd69}:		p = 14'd345;
            {7'd5,7'd70}:		p = 14'd350;
            {7'd5,7'd71}:		p = 14'd355;
            {7'd5,7'd72}:		p = 14'd360;
            {7'd5,7'd73}:		p = 14'd365;
            {7'd5,7'd74}:		p = 14'd370;
            {7'd5,7'd75}:		p = 14'd375;
            {7'd5,7'd76}:		p = 14'd380;
            {7'd5,7'd77}:		p = 14'd385;
            {7'd5,7'd78}:		p = 14'd390;
            {7'd5,7'd79}:		p = 14'd395;
            {7'd5,7'd80}:		p = 14'd400;
            {7'd5,7'd81}:		p = 14'd405;
            {7'd5,7'd82}:		p = 14'd410;
            {7'd5,7'd83}:		p = 14'd415;
            {7'd5,7'd84}:		p = 14'd420;
            {7'd5,7'd85}:		p = 14'd425;
            {7'd5,7'd86}:		p = 14'd430;
            {7'd5,7'd87}:		p = 14'd435;
            {7'd5,7'd88}:		p = 14'd440;
            {7'd5,7'd89}:		p = 14'd445;
            {7'd5,7'd90}:		p = 14'd450;
            {7'd5,7'd91}:		p = 14'd455;
            {7'd5,7'd92}:		p = 14'd460;
            {7'd5,7'd93}:		p = 14'd465;
            {7'd5,7'd94}:		p = 14'd470;
            {7'd5,7'd95}:		p = 14'd475;
            {7'd5,7'd96}:		p = 14'd480;
            {7'd5,7'd97}:		p = 14'd485;
            {7'd5,7'd98}:		p = 14'd490;
            {7'd5,7'd99}:		p = 14'd495;
            {7'd5,7'd100}:		p = 14'd500;
            {7'd5,7'd101}:		p = 14'd505;
            {7'd5,7'd102}:		p = 14'd510;
            {7'd5,7'd103}:		p = 14'd515;
            {7'd5,7'd104}:		p = 14'd520;
            {7'd5,7'd105}:		p = 14'd525;
            {7'd5,7'd106}:		p = 14'd530;
            {7'd5,7'd107}:		p = 14'd535;
            {7'd5,7'd108}:		p = 14'd540;
            {7'd5,7'd109}:		p = 14'd545;
            {7'd5,7'd110}:		p = 14'd550;
            {7'd5,7'd111}:		p = 14'd555;
            {7'd5,7'd112}:		p = 14'd560;
            {7'd5,7'd113}:		p = 14'd565;
            {7'd5,7'd114}:		p = 14'd570;
            {7'd5,7'd115}:		p = 14'd575;
            {7'd5,7'd116}:		p = 14'd580;
            {7'd5,7'd117}:		p = 14'd585;
            {7'd5,7'd118}:		p = 14'd590;
            {7'd5,7'd119}:		p = 14'd595;
            {7'd5,7'd120}:		p = 14'd600;
            {7'd5,7'd121}:		p = 14'd605;
            {7'd5,7'd122}:		p = 14'd610;
            {7'd5,7'd123}:		p = 14'd615;
            {7'd5,7'd124}:		p = 14'd620;
            {7'd5,7'd125}:		p = 14'd625;
            {7'd5,7'd126}:		p = 14'd630;
            {7'd5,7'd127}:		p = 14'd635;
            {7'd6,7'd0}:		p = 14'd0;
            {7'd6,7'd1}:		p = 14'd6;
            {7'd6,7'd2}:		p = 14'd12;
            {7'd6,7'd3}:		p = 14'd18;
            {7'd6,7'd4}:		p = 14'd24;
            {7'd6,7'd5}:		p = 14'd30;
            {7'd6,7'd6}:		p = 14'd36;
            {7'd6,7'd7}:		p = 14'd42;
            {7'd6,7'd8}:		p = 14'd48;
            {7'd6,7'd9}:		p = 14'd54;
            {7'd6,7'd10}:		p = 14'd60;
            {7'd6,7'd11}:		p = 14'd66;
            {7'd6,7'd12}:		p = 14'd72;
            {7'd6,7'd13}:		p = 14'd78;
            {7'd6,7'd14}:		p = 14'd84;
            {7'd6,7'd15}:		p = 14'd90;
            {7'd6,7'd16}:		p = 14'd96;
            {7'd6,7'd17}:		p = 14'd102;
            {7'd6,7'd18}:		p = 14'd108;
            {7'd6,7'd19}:		p = 14'd114;
            {7'd6,7'd20}:		p = 14'd120;
            {7'd6,7'd21}:		p = 14'd126;
            {7'd6,7'd22}:		p = 14'd132;
            {7'd6,7'd23}:		p = 14'd138;
            {7'd6,7'd24}:		p = 14'd144;
            {7'd6,7'd25}:		p = 14'd150;
            {7'd6,7'd26}:		p = 14'd156;
            {7'd6,7'd27}:		p = 14'd162;
            {7'd6,7'd28}:		p = 14'd168;
            {7'd6,7'd29}:		p = 14'd174;
            {7'd6,7'd30}:		p = 14'd180;
            {7'd6,7'd31}:		p = 14'd186;
            {7'd6,7'd32}:		p = 14'd192;
            {7'd6,7'd33}:		p = 14'd198;
            {7'd6,7'd34}:		p = 14'd204;
            {7'd6,7'd35}:		p = 14'd210;
            {7'd6,7'd36}:		p = 14'd216;
            {7'd6,7'd37}:		p = 14'd222;
            {7'd6,7'd38}:		p = 14'd228;
            {7'd6,7'd39}:		p = 14'd234;
            {7'd6,7'd40}:		p = 14'd240;
            {7'd6,7'd41}:		p = 14'd246;
            {7'd6,7'd42}:		p = 14'd252;
            {7'd6,7'd43}:		p = 14'd258;
            {7'd6,7'd44}:		p = 14'd264;
            {7'd6,7'd45}:		p = 14'd270;
            {7'd6,7'd46}:		p = 14'd276;
            {7'd6,7'd47}:		p = 14'd282;
            {7'd6,7'd48}:		p = 14'd288;
            {7'd6,7'd49}:		p = 14'd294;
            {7'd6,7'd50}:		p = 14'd300;
            {7'd6,7'd51}:		p = 14'd306;
            {7'd6,7'd52}:		p = 14'd312;
            {7'd6,7'd53}:		p = 14'd318;
            {7'd6,7'd54}:		p = 14'd324;
            {7'd6,7'd55}:		p = 14'd330;
            {7'd6,7'd56}:		p = 14'd336;
            {7'd6,7'd57}:		p = 14'd342;
            {7'd6,7'd58}:		p = 14'd348;
            {7'd6,7'd59}:		p = 14'd354;
            {7'd6,7'd60}:		p = 14'd360;
            {7'd6,7'd61}:		p = 14'd366;
            {7'd6,7'd62}:		p = 14'd372;
            {7'd6,7'd63}:		p = 14'd378;
            {7'd6,7'd64}:		p = 14'd384;
            {7'd6,7'd65}:		p = 14'd390;
            {7'd6,7'd66}:		p = 14'd396;
            {7'd6,7'd67}:		p = 14'd402;
            {7'd6,7'd68}:		p = 14'd408;
            {7'd6,7'd69}:		p = 14'd414;
            {7'd6,7'd70}:		p = 14'd420;
            {7'd6,7'd71}:		p = 14'd426;
            {7'd6,7'd72}:		p = 14'd432;
            {7'd6,7'd73}:		p = 14'd438;
            {7'd6,7'd74}:		p = 14'd444;
            {7'd6,7'd75}:		p = 14'd450;
            {7'd6,7'd76}:		p = 14'd456;
            {7'd6,7'd77}:		p = 14'd462;
            {7'd6,7'd78}:		p = 14'd468;
            {7'd6,7'd79}:		p = 14'd474;
            {7'd6,7'd80}:		p = 14'd480;
            {7'd6,7'd81}:		p = 14'd486;
            {7'd6,7'd82}:		p = 14'd492;
            {7'd6,7'd83}:		p = 14'd498;
            {7'd6,7'd84}:		p = 14'd504;
            {7'd6,7'd85}:		p = 14'd510;
            {7'd6,7'd86}:		p = 14'd516;
            {7'd6,7'd87}:		p = 14'd522;
            {7'd6,7'd88}:		p = 14'd528;
            {7'd6,7'd89}:		p = 14'd534;
            {7'd6,7'd90}:		p = 14'd540;
            {7'd6,7'd91}:		p = 14'd546;
            {7'd6,7'd92}:		p = 14'd552;
            {7'd6,7'd93}:		p = 14'd558;
            {7'd6,7'd94}:		p = 14'd564;
            {7'd6,7'd95}:		p = 14'd570;
            {7'd6,7'd96}:		p = 14'd576;
            {7'd6,7'd97}:		p = 14'd582;
            {7'd6,7'd98}:		p = 14'd588;
            {7'd6,7'd99}:		p = 14'd594;
            {7'd6,7'd100}:		p = 14'd600;
            {7'd6,7'd101}:		p = 14'd606;
            {7'd6,7'd102}:		p = 14'd612;
            {7'd6,7'd103}:		p = 14'd618;
            {7'd6,7'd104}:		p = 14'd624;
            {7'd6,7'd105}:		p = 14'd630;
            {7'd6,7'd106}:		p = 14'd636;
            {7'd6,7'd107}:		p = 14'd642;
            {7'd6,7'd108}:		p = 14'd648;
            {7'd6,7'd109}:		p = 14'd654;
            {7'd6,7'd110}:		p = 14'd660;
            {7'd6,7'd111}:		p = 14'd666;
            {7'd6,7'd112}:		p = 14'd672;
            {7'd6,7'd113}:		p = 14'd678;
            {7'd6,7'd114}:		p = 14'd684;
            {7'd6,7'd115}:		p = 14'd690;
            {7'd6,7'd116}:		p = 14'd696;
            {7'd6,7'd117}:		p = 14'd702;
            {7'd6,7'd118}:		p = 14'd708;
            {7'd6,7'd119}:		p = 14'd714;
            {7'd6,7'd120}:		p = 14'd720;
            {7'd6,7'd121}:		p = 14'd726;
            {7'd6,7'd122}:		p = 14'd732;
            {7'd6,7'd123}:		p = 14'd738;
            {7'd6,7'd124}:		p = 14'd744;
            {7'd6,7'd125}:		p = 14'd750;
            {7'd6,7'd126}:		p = 14'd756;
            {7'd6,7'd127}:		p = 14'd762;
            {7'd7,7'd0}:		p = 14'd0;
            {7'd7,7'd1}:		p = 14'd7;
            {7'd7,7'd2}:		p = 14'd14;
            {7'd7,7'd3}:		p = 14'd21;
            {7'd7,7'd4}:		p = 14'd28;
            {7'd7,7'd5}:		p = 14'd35;
            {7'd7,7'd6}:		p = 14'd42;
            {7'd7,7'd7}:		p = 14'd49;
            {7'd7,7'd8}:		p = 14'd56;
            {7'd7,7'd9}:		p = 14'd63;
            {7'd7,7'd10}:		p = 14'd70;
            {7'd7,7'd11}:		p = 14'd77;
            {7'd7,7'd12}:		p = 14'd84;
            {7'd7,7'd13}:		p = 14'd91;
            {7'd7,7'd14}:		p = 14'd98;
            {7'd7,7'd15}:		p = 14'd105;
            {7'd7,7'd16}:		p = 14'd112;
            {7'd7,7'd17}:		p = 14'd119;
            {7'd7,7'd18}:		p = 14'd126;
            {7'd7,7'd19}:		p = 14'd133;
            {7'd7,7'd20}:		p = 14'd140;
            {7'd7,7'd21}:		p = 14'd147;
            {7'd7,7'd22}:		p = 14'd154;
            {7'd7,7'd23}:		p = 14'd161;
            {7'd7,7'd24}:		p = 14'd168;
            {7'd7,7'd25}:		p = 14'd175;
            {7'd7,7'd26}:		p = 14'd182;
            {7'd7,7'd27}:		p = 14'd189;
            {7'd7,7'd28}:		p = 14'd196;
            {7'd7,7'd29}:		p = 14'd203;
            {7'd7,7'd30}:		p = 14'd210;
            {7'd7,7'd31}:		p = 14'd217;
            {7'd7,7'd32}:		p = 14'd224;
            {7'd7,7'd33}:		p = 14'd231;
            {7'd7,7'd34}:		p = 14'd238;
            {7'd7,7'd35}:		p = 14'd245;
            {7'd7,7'd36}:		p = 14'd252;
            {7'd7,7'd37}:		p = 14'd259;
            {7'd7,7'd38}:		p = 14'd266;
            {7'd7,7'd39}:		p = 14'd273;
            {7'd7,7'd40}:		p = 14'd280;
            {7'd7,7'd41}:		p = 14'd287;
            {7'd7,7'd42}:		p = 14'd294;
            {7'd7,7'd43}:		p = 14'd301;
            {7'd7,7'd44}:		p = 14'd308;
            {7'd7,7'd45}:		p = 14'd315;
            {7'd7,7'd46}:		p = 14'd322;
            {7'd7,7'd47}:		p = 14'd329;
            {7'd7,7'd48}:		p = 14'd336;
            {7'd7,7'd49}:		p = 14'd343;
            {7'd7,7'd50}:		p = 14'd350;
            {7'd7,7'd51}:		p = 14'd357;
            {7'd7,7'd52}:		p = 14'd364;
            {7'd7,7'd53}:		p = 14'd371;
            {7'd7,7'd54}:		p = 14'd378;
            {7'd7,7'd55}:		p = 14'd385;
            {7'd7,7'd56}:		p = 14'd392;
            {7'd7,7'd57}:		p = 14'd399;
            {7'd7,7'd58}:		p = 14'd406;
            {7'd7,7'd59}:		p = 14'd413;
            {7'd7,7'd60}:		p = 14'd420;
            {7'd7,7'd61}:		p = 14'd427;
            {7'd7,7'd62}:		p = 14'd434;
            {7'd7,7'd63}:		p = 14'd441;
            {7'd7,7'd64}:		p = 14'd448;
            {7'd7,7'd65}:		p = 14'd455;
            {7'd7,7'd66}:		p = 14'd462;
            {7'd7,7'd67}:		p = 14'd469;
            {7'd7,7'd68}:		p = 14'd476;
            {7'd7,7'd69}:		p = 14'd483;
            {7'd7,7'd70}:		p = 14'd490;
            {7'd7,7'd71}:		p = 14'd497;
            {7'd7,7'd72}:		p = 14'd504;
            {7'd7,7'd73}:		p = 14'd511;
            {7'd7,7'd74}:		p = 14'd518;
            {7'd7,7'd75}:		p = 14'd525;
            {7'd7,7'd76}:		p = 14'd532;
            {7'd7,7'd77}:		p = 14'd539;
            {7'd7,7'd78}:		p = 14'd546;
            {7'd7,7'd79}:		p = 14'd553;
            {7'd7,7'd80}:		p = 14'd560;
            {7'd7,7'd81}:		p = 14'd567;
            {7'd7,7'd82}:		p = 14'd574;
            {7'd7,7'd83}:		p = 14'd581;
            {7'd7,7'd84}:		p = 14'd588;
            {7'd7,7'd85}:		p = 14'd595;
            {7'd7,7'd86}:		p = 14'd602;
            {7'd7,7'd87}:		p = 14'd609;
            {7'd7,7'd88}:		p = 14'd616;
            {7'd7,7'd89}:		p = 14'd623;
            {7'd7,7'd90}:		p = 14'd630;
            {7'd7,7'd91}:		p = 14'd637;
            {7'd7,7'd92}:		p = 14'd644;
            {7'd7,7'd93}:		p = 14'd651;
            {7'd7,7'd94}:		p = 14'd658;
            {7'd7,7'd95}:		p = 14'd665;
            {7'd7,7'd96}:		p = 14'd672;
            {7'd7,7'd97}:		p = 14'd679;
            {7'd7,7'd98}:		p = 14'd686;
            {7'd7,7'd99}:		p = 14'd693;
            {7'd7,7'd100}:		p = 14'd700;
            {7'd7,7'd101}:		p = 14'd707;
            {7'd7,7'd102}:		p = 14'd714;
            {7'd7,7'd103}:		p = 14'd721;
            {7'd7,7'd104}:		p = 14'd728;
            {7'd7,7'd105}:		p = 14'd735;
            {7'd7,7'd106}:		p = 14'd742;
            {7'd7,7'd107}:		p = 14'd749;
            {7'd7,7'd108}:		p = 14'd756;
            {7'd7,7'd109}:		p = 14'd763;
            {7'd7,7'd110}:		p = 14'd770;
            {7'd7,7'd111}:		p = 14'd777;
            {7'd7,7'd112}:		p = 14'd784;
            {7'd7,7'd113}:		p = 14'd791;
            {7'd7,7'd114}:		p = 14'd798;
            {7'd7,7'd115}:		p = 14'd805;
            {7'd7,7'd116}:		p = 14'd812;
            {7'd7,7'd117}:		p = 14'd819;
            {7'd7,7'd118}:		p = 14'd826;
            {7'd7,7'd119}:		p = 14'd833;
            {7'd7,7'd120}:		p = 14'd840;
            {7'd7,7'd121}:		p = 14'd847;
            {7'd7,7'd122}:		p = 14'd854;
            {7'd7,7'd123}:		p = 14'd861;
            {7'd7,7'd124}:		p = 14'd868;
            {7'd7,7'd125}:		p = 14'd875;
            {7'd7,7'd126}:		p = 14'd882;
            {7'd7,7'd127}:		p = 14'd889;
            {7'd8,7'd0}:		p = 14'd0;
            {7'd8,7'd1}:		p = 14'd8;
            {7'd8,7'd2}:		p = 14'd16;
            {7'd8,7'd3}:		p = 14'd24;
            {7'd8,7'd4}:		p = 14'd32;
            {7'd8,7'd5}:		p = 14'd40;
            {7'd8,7'd6}:		p = 14'd48;
            {7'd8,7'd7}:		p = 14'd56;
            {7'd8,7'd8}:		p = 14'd64;
            {7'd8,7'd9}:		p = 14'd72;
            {7'd8,7'd10}:		p = 14'd80;
            {7'd8,7'd11}:		p = 14'd88;
            {7'd8,7'd12}:		p = 14'd96;
            {7'd8,7'd13}:		p = 14'd104;
            {7'd8,7'd14}:		p = 14'd112;
            {7'd8,7'd15}:		p = 14'd120;
            {7'd8,7'd16}:		p = 14'd128;
            {7'd8,7'd17}:		p = 14'd136;
            {7'd8,7'd18}:		p = 14'd144;
            {7'd8,7'd19}:		p = 14'd152;
            {7'd8,7'd20}:		p = 14'd160;
            {7'd8,7'd21}:		p = 14'd168;
            {7'd8,7'd22}:		p = 14'd176;
            {7'd8,7'd23}:		p = 14'd184;
            {7'd8,7'd24}:		p = 14'd192;
            {7'd8,7'd25}:		p = 14'd200;
            {7'd8,7'd26}:		p = 14'd208;
            {7'd8,7'd27}:		p = 14'd216;
            {7'd8,7'd28}:		p = 14'd224;
            {7'd8,7'd29}:		p = 14'd232;
            {7'd8,7'd30}:		p = 14'd240;
            {7'd8,7'd31}:		p = 14'd248;
            {7'd8,7'd32}:		p = 14'd256;
            {7'd8,7'd33}:		p = 14'd264;
            {7'd8,7'd34}:		p = 14'd272;
            {7'd8,7'd35}:		p = 14'd280;
            {7'd8,7'd36}:		p = 14'd288;
            {7'd8,7'd37}:		p = 14'd296;
            {7'd8,7'd38}:		p = 14'd304;
            {7'd8,7'd39}:		p = 14'd312;
            {7'd8,7'd40}:		p = 14'd320;
            {7'd8,7'd41}:		p = 14'd328;
            {7'd8,7'd42}:		p = 14'd336;
            {7'd8,7'd43}:		p = 14'd344;
            {7'd8,7'd44}:		p = 14'd352;
            {7'd8,7'd45}:		p = 14'd360;
            {7'd8,7'd46}:		p = 14'd368;
            {7'd8,7'd47}:		p = 14'd376;
            {7'd8,7'd48}:		p = 14'd384;
            {7'd8,7'd49}:		p = 14'd392;
            {7'd8,7'd50}:		p = 14'd400;
            {7'd8,7'd51}:		p = 14'd408;
            {7'd8,7'd52}:		p = 14'd416;
            {7'd8,7'd53}:		p = 14'd424;
            {7'd8,7'd54}:		p = 14'd432;
            {7'd8,7'd55}:		p = 14'd440;
            {7'd8,7'd56}:		p = 14'd448;
            {7'd8,7'd57}:		p = 14'd456;
            {7'd8,7'd58}:		p = 14'd464;
            {7'd8,7'd59}:		p = 14'd472;
            {7'd8,7'd60}:		p = 14'd480;
            {7'd8,7'd61}:		p = 14'd488;
            {7'd8,7'd62}:		p = 14'd496;
            {7'd8,7'd63}:		p = 14'd504;
            {7'd8,7'd64}:		p = 14'd512;
            {7'd8,7'd65}:		p = 14'd520;
            {7'd8,7'd66}:		p = 14'd528;
            {7'd8,7'd67}:		p = 14'd536;
            {7'd8,7'd68}:		p = 14'd544;
            {7'd8,7'd69}:		p = 14'd552;
            {7'd8,7'd70}:		p = 14'd560;
            {7'd8,7'd71}:		p = 14'd568;
            {7'd8,7'd72}:		p = 14'd576;
            {7'd8,7'd73}:		p = 14'd584;
            {7'd8,7'd74}:		p = 14'd592;
            {7'd8,7'd75}:		p = 14'd600;
            {7'd8,7'd76}:		p = 14'd608;
            {7'd8,7'd77}:		p = 14'd616;
            {7'd8,7'd78}:		p = 14'd624;
            {7'd8,7'd79}:		p = 14'd632;
            {7'd8,7'd80}:		p = 14'd640;
            {7'd8,7'd81}:		p = 14'd648;
            {7'd8,7'd82}:		p = 14'd656;
            {7'd8,7'd83}:		p = 14'd664;
            {7'd8,7'd84}:		p = 14'd672;
            {7'd8,7'd85}:		p = 14'd680;
            {7'd8,7'd86}:		p = 14'd688;
            {7'd8,7'd87}:		p = 14'd696;
            {7'd8,7'd88}:		p = 14'd704;
            {7'd8,7'd89}:		p = 14'd712;
            {7'd8,7'd90}:		p = 14'd720;
            {7'd8,7'd91}:		p = 14'd728;
            {7'd8,7'd92}:		p = 14'd736;
            {7'd8,7'd93}:		p = 14'd744;
            {7'd8,7'd94}:		p = 14'd752;
            {7'd8,7'd95}:		p = 14'd760;
            {7'd8,7'd96}:		p = 14'd768;
            {7'd8,7'd97}:		p = 14'd776;
            {7'd8,7'd98}:		p = 14'd784;
            {7'd8,7'd99}:		p = 14'd792;
            {7'd8,7'd100}:		p = 14'd800;
            {7'd8,7'd101}:		p = 14'd808;
            {7'd8,7'd102}:		p = 14'd816;
            {7'd8,7'd103}:		p = 14'd824;
            {7'd8,7'd104}:		p = 14'd832;
            {7'd8,7'd105}:		p = 14'd840;
            {7'd8,7'd106}:		p = 14'd848;
            {7'd8,7'd107}:		p = 14'd856;
            {7'd8,7'd108}:		p = 14'd864;
            {7'd8,7'd109}:		p = 14'd872;
            {7'd8,7'd110}:		p = 14'd880;
            {7'd8,7'd111}:		p = 14'd888;
            {7'd8,7'd112}:		p = 14'd896;
            {7'd8,7'd113}:		p = 14'd904;
            {7'd8,7'd114}:		p = 14'd912;
            {7'd8,7'd115}:		p = 14'd920;
            {7'd8,7'd116}:		p = 14'd928;
            {7'd8,7'd117}:		p = 14'd936;
            {7'd8,7'd118}:		p = 14'd944;
            {7'd8,7'd119}:		p = 14'd952;
            {7'd8,7'd120}:		p = 14'd960;
            {7'd8,7'd121}:		p = 14'd968;
            {7'd8,7'd122}:		p = 14'd976;
            {7'd8,7'd123}:		p = 14'd984;
            {7'd8,7'd124}:		p = 14'd992;
            {7'd8,7'd125}:		p = 14'd1000;
            {7'd8,7'd126}:		p = 14'd1008;
            {7'd8,7'd127}:		p = 14'd1016;
            {7'd9,7'd0}:		p = 14'd0;
            {7'd9,7'd1}:		p = 14'd9;
            {7'd9,7'd2}:		p = 14'd18;
            {7'd9,7'd3}:		p = 14'd27;
            {7'd9,7'd4}:		p = 14'd36;
            {7'd9,7'd5}:		p = 14'd45;
            {7'd9,7'd6}:		p = 14'd54;
            {7'd9,7'd7}:		p = 14'd63;
            {7'd9,7'd8}:		p = 14'd72;
            {7'd9,7'd9}:		p = 14'd81;
            {7'd9,7'd10}:		p = 14'd90;
            {7'd9,7'd11}:		p = 14'd99;
            {7'd9,7'd12}:		p = 14'd108;
            {7'd9,7'd13}:		p = 14'd117;
            {7'd9,7'd14}:		p = 14'd126;
            {7'd9,7'd15}:		p = 14'd135;
            {7'd9,7'd16}:		p = 14'd144;
            {7'd9,7'd17}:		p = 14'd153;
            {7'd9,7'd18}:		p = 14'd162;
            {7'd9,7'd19}:		p = 14'd171;
            {7'd9,7'd20}:		p = 14'd180;
            {7'd9,7'd21}:		p = 14'd189;
            {7'd9,7'd22}:		p = 14'd198;
            {7'd9,7'd23}:		p = 14'd207;
            {7'd9,7'd24}:		p = 14'd216;
            {7'd9,7'd25}:		p = 14'd225;
            {7'd9,7'd26}:		p = 14'd234;
            {7'd9,7'd27}:		p = 14'd243;
            {7'd9,7'd28}:		p = 14'd252;
            {7'd9,7'd29}:		p = 14'd261;
            {7'd9,7'd30}:		p = 14'd270;
            {7'd9,7'd31}:		p = 14'd279;
            {7'd9,7'd32}:		p = 14'd288;
            {7'd9,7'd33}:		p = 14'd297;
            {7'd9,7'd34}:		p = 14'd306;
            {7'd9,7'd35}:		p = 14'd315;
            {7'd9,7'd36}:		p = 14'd324;
            {7'd9,7'd37}:		p = 14'd333;
            {7'd9,7'd38}:		p = 14'd342;
            {7'd9,7'd39}:		p = 14'd351;
            {7'd9,7'd40}:		p = 14'd360;
            {7'd9,7'd41}:		p = 14'd369;
            {7'd9,7'd42}:		p = 14'd378;
            {7'd9,7'd43}:		p = 14'd387;
            {7'd9,7'd44}:		p = 14'd396;
            {7'd9,7'd45}:		p = 14'd405;
            {7'd9,7'd46}:		p = 14'd414;
            {7'd9,7'd47}:		p = 14'd423;
            {7'd9,7'd48}:		p = 14'd432;
            {7'd9,7'd49}:		p = 14'd441;
            {7'd9,7'd50}:		p = 14'd450;
            {7'd9,7'd51}:		p = 14'd459;
            {7'd9,7'd52}:		p = 14'd468;
            {7'd9,7'd53}:		p = 14'd477;
            {7'd9,7'd54}:		p = 14'd486;
            {7'd9,7'd55}:		p = 14'd495;
            {7'd9,7'd56}:		p = 14'd504;
            {7'd9,7'd57}:		p = 14'd513;
            {7'd9,7'd58}:		p = 14'd522;
            {7'd9,7'd59}:		p = 14'd531;
            {7'd9,7'd60}:		p = 14'd540;
            {7'd9,7'd61}:		p = 14'd549;
            {7'd9,7'd62}:		p = 14'd558;
            {7'd9,7'd63}:		p = 14'd567;
            {7'd9,7'd64}:		p = 14'd576;
            {7'd9,7'd65}:		p = 14'd585;
            {7'd9,7'd66}:		p = 14'd594;
            {7'd9,7'd67}:		p = 14'd603;
            {7'd9,7'd68}:		p = 14'd612;
            {7'd9,7'd69}:		p = 14'd621;
            {7'd9,7'd70}:		p = 14'd630;
            {7'd9,7'd71}:		p = 14'd639;
            {7'd9,7'd72}:		p = 14'd648;
            {7'd9,7'd73}:		p = 14'd657;
            {7'd9,7'd74}:		p = 14'd666;
            {7'd9,7'd75}:		p = 14'd675;
            {7'd9,7'd76}:		p = 14'd684;
            {7'd9,7'd77}:		p = 14'd693;
            {7'd9,7'd78}:		p = 14'd702;
            {7'd9,7'd79}:		p = 14'd711;
            {7'd9,7'd80}:		p = 14'd720;
            {7'd9,7'd81}:		p = 14'd729;
            {7'd9,7'd82}:		p = 14'd738;
            {7'd9,7'd83}:		p = 14'd747;
            {7'd9,7'd84}:		p = 14'd756;
            {7'd9,7'd85}:		p = 14'd765;
            {7'd9,7'd86}:		p = 14'd774;
            {7'd9,7'd87}:		p = 14'd783;
            {7'd9,7'd88}:		p = 14'd792;
            {7'd9,7'd89}:		p = 14'd801;
            {7'd9,7'd90}:		p = 14'd810;
            {7'd9,7'd91}:		p = 14'd819;
            {7'd9,7'd92}:		p = 14'd828;
            {7'd9,7'd93}:		p = 14'd837;
            {7'd9,7'd94}:		p = 14'd846;
            {7'd9,7'd95}:		p = 14'd855;
            {7'd9,7'd96}:		p = 14'd864;
            {7'd9,7'd97}:		p = 14'd873;
            {7'd9,7'd98}:		p = 14'd882;
            {7'd9,7'd99}:		p = 14'd891;
            {7'd9,7'd100}:		p = 14'd900;
            {7'd9,7'd101}:		p = 14'd909;
            {7'd9,7'd102}:		p = 14'd918;
            {7'd9,7'd103}:		p = 14'd927;
            {7'd9,7'd104}:		p = 14'd936;
            {7'd9,7'd105}:		p = 14'd945;
            {7'd9,7'd106}:		p = 14'd954;
            {7'd9,7'd107}:		p = 14'd963;
            {7'd9,7'd108}:		p = 14'd972;
            {7'd9,7'd109}:		p = 14'd981;
            {7'd9,7'd110}:		p = 14'd990;
            {7'd9,7'd111}:		p = 14'd999;
            {7'd9,7'd112}:		p = 14'd1008;
            {7'd9,7'd113}:		p = 14'd1017;
            {7'd9,7'd114}:		p = 14'd1026;
            {7'd9,7'd115}:		p = 14'd1035;
            {7'd9,7'd116}:		p = 14'd1044;
            {7'd9,7'd117}:		p = 14'd1053;
            {7'd9,7'd118}:		p = 14'd1062;
            {7'd9,7'd119}:		p = 14'd1071;
            {7'd9,7'd120}:		p = 14'd1080;
            {7'd9,7'd121}:		p = 14'd1089;
            {7'd9,7'd122}:		p = 14'd1098;
            {7'd9,7'd123}:		p = 14'd1107;
            {7'd9,7'd124}:		p = 14'd1116;
            {7'd9,7'd125}:		p = 14'd1125;
            {7'd9,7'd126}:		p = 14'd1134;
            {7'd9,7'd127}:		p = 14'd1143;
            {7'd10,7'd0}:		p = 14'd0;
            {7'd10,7'd1}:		p = 14'd10;
            {7'd10,7'd2}:		p = 14'd20;
            {7'd10,7'd3}:		p = 14'd30;
            {7'd10,7'd4}:		p = 14'd40;
            {7'd10,7'd5}:		p = 14'd50;
            {7'd10,7'd6}:		p = 14'd60;
            {7'd10,7'd7}:		p = 14'd70;
            {7'd10,7'd8}:		p = 14'd80;
            {7'd10,7'd9}:		p = 14'd90;
            {7'd10,7'd10}:		p = 14'd100;
            {7'd10,7'd11}:		p = 14'd110;
            {7'd10,7'd12}:		p = 14'd120;
            {7'd10,7'd13}:		p = 14'd130;
            {7'd10,7'd14}:		p = 14'd140;
            {7'd10,7'd15}:		p = 14'd150;
            {7'd10,7'd16}:		p = 14'd160;
            {7'd10,7'd17}:		p = 14'd170;
            {7'd10,7'd18}:		p = 14'd180;
            {7'd10,7'd19}:		p = 14'd190;
            {7'd10,7'd20}:		p = 14'd200;
            {7'd10,7'd21}:		p = 14'd210;
            {7'd10,7'd22}:		p = 14'd220;
            {7'd10,7'd23}:		p = 14'd230;
            {7'd10,7'd24}:		p = 14'd240;
            {7'd10,7'd25}:		p = 14'd250;
            {7'd10,7'd26}:		p = 14'd260;
            {7'd10,7'd27}:		p = 14'd270;
            {7'd10,7'd28}:		p = 14'd280;
            {7'd10,7'd29}:		p = 14'd290;
            {7'd10,7'd30}:		p = 14'd300;
            {7'd10,7'd31}:		p = 14'd310;
            {7'd10,7'd32}:		p = 14'd320;
            {7'd10,7'd33}:		p = 14'd330;
            {7'd10,7'd34}:		p = 14'd340;
            {7'd10,7'd35}:		p = 14'd350;
            {7'd10,7'd36}:		p = 14'd360;
            {7'd10,7'd37}:		p = 14'd370;
            {7'd10,7'd38}:		p = 14'd380;
            {7'd10,7'd39}:		p = 14'd390;
            {7'd10,7'd40}:		p = 14'd400;
            {7'd10,7'd41}:		p = 14'd410;
            {7'd10,7'd42}:		p = 14'd420;
            {7'd10,7'd43}:		p = 14'd430;
            {7'd10,7'd44}:		p = 14'd440;
            {7'd10,7'd45}:		p = 14'd450;
            {7'd10,7'd46}:		p = 14'd460;
            {7'd10,7'd47}:		p = 14'd470;
            {7'd10,7'd48}:		p = 14'd480;
            {7'd10,7'd49}:		p = 14'd490;
            {7'd10,7'd50}:		p = 14'd500;
            {7'd10,7'd51}:		p = 14'd510;
            {7'd10,7'd52}:		p = 14'd520;
            {7'd10,7'd53}:		p = 14'd530;
            {7'd10,7'd54}:		p = 14'd540;
            {7'd10,7'd55}:		p = 14'd550;
            {7'd10,7'd56}:		p = 14'd560;
            {7'd10,7'd57}:		p = 14'd570;
            {7'd10,7'd58}:		p = 14'd580;
            {7'd10,7'd59}:		p = 14'd590;
            {7'd10,7'd60}:		p = 14'd600;
            {7'd10,7'd61}:		p = 14'd610;
            {7'd10,7'd62}:		p = 14'd620;
            {7'd10,7'd63}:		p = 14'd630;
            {7'd10,7'd64}:		p = 14'd640;
            {7'd10,7'd65}:		p = 14'd650;
            {7'd10,7'd66}:		p = 14'd660;
            {7'd10,7'd67}:		p = 14'd670;
            {7'd10,7'd68}:		p = 14'd680;
            {7'd10,7'd69}:		p = 14'd690;
            {7'd10,7'd70}:		p = 14'd700;
            {7'd10,7'd71}:		p = 14'd710;
            {7'd10,7'd72}:		p = 14'd720;
            {7'd10,7'd73}:		p = 14'd730;
            {7'd10,7'd74}:		p = 14'd740;
            {7'd10,7'd75}:		p = 14'd750;
            {7'd10,7'd76}:		p = 14'd760;
            {7'd10,7'd77}:		p = 14'd770;
            {7'd10,7'd78}:		p = 14'd780;
            {7'd10,7'd79}:		p = 14'd790;
            {7'd10,7'd80}:		p = 14'd800;
            {7'd10,7'd81}:		p = 14'd810;
            {7'd10,7'd82}:		p = 14'd820;
            {7'd10,7'd83}:		p = 14'd830;
            {7'd10,7'd84}:		p = 14'd840;
            {7'd10,7'd85}:		p = 14'd850;
            {7'd10,7'd86}:		p = 14'd860;
            {7'd10,7'd87}:		p = 14'd870;
            {7'd10,7'd88}:		p = 14'd880;
            {7'd10,7'd89}:		p = 14'd890;
            {7'd10,7'd90}:		p = 14'd900;
            {7'd10,7'd91}:		p = 14'd910;
            {7'd10,7'd92}:		p = 14'd920;
            {7'd10,7'd93}:		p = 14'd930;
            {7'd10,7'd94}:		p = 14'd940;
            {7'd10,7'd95}:		p = 14'd950;
            {7'd10,7'd96}:		p = 14'd960;
            {7'd10,7'd97}:		p = 14'd970;
            {7'd10,7'd98}:		p = 14'd980;
            {7'd10,7'd99}:		p = 14'd990;
            {7'd10,7'd100}:		p = 14'd1000;
            {7'd10,7'd101}:		p = 14'd1010;
            {7'd10,7'd102}:		p = 14'd1020;
            {7'd10,7'd103}:		p = 14'd1030;
            {7'd10,7'd104}:		p = 14'd1040;
            {7'd10,7'd105}:		p = 14'd1050;
            {7'd10,7'd106}:		p = 14'd1060;
            {7'd10,7'd107}:		p = 14'd1070;
            {7'd10,7'd108}:		p = 14'd1080;
            {7'd10,7'd109}:		p = 14'd1090;
            {7'd10,7'd110}:		p = 14'd1100;
            {7'd10,7'd111}:		p = 14'd1110;
            {7'd10,7'd112}:		p = 14'd1120;
            {7'd10,7'd113}:		p = 14'd1130;
            {7'd10,7'd114}:		p = 14'd1140;
            {7'd10,7'd115}:		p = 14'd1150;
            {7'd10,7'd116}:		p = 14'd1160;
            {7'd10,7'd117}:		p = 14'd1170;
            {7'd10,7'd118}:		p = 14'd1180;
            {7'd10,7'd119}:		p = 14'd1190;
            {7'd10,7'd120}:		p = 14'd1200;
            {7'd10,7'd121}:		p = 14'd1210;
            {7'd10,7'd122}:		p = 14'd1220;
            {7'd10,7'd123}:		p = 14'd1230;
            {7'd10,7'd124}:		p = 14'd1240;
            {7'd10,7'd125}:		p = 14'd1250;
            {7'd10,7'd126}:		p = 14'd1260;
            {7'd10,7'd127}:		p = 14'd1270;
            {7'd11,7'd0}:		p = 14'd0;
            {7'd11,7'd1}:		p = 14'd11;
            {7'd11,7'd2}:		p = 14'd22;
            {7'd11,7'd3}:		p = 14'd33;
            {7'd11,7'd4}:		p = 14'd44;
            {7'd11,7'd5}:		p = 14'd55;
            {7'd11,7'd6}:		p = 14'd66;
            {7'd11,7'd7}:		p = 14'd77;
            {7'd11,7'd8}:		p = 14'd88;
            {7'd11,7'd9}:		p = 14'd99;
            {7'd11,7'd10}:		p = 14'd110;
            {7'd11,7'd11}:		p = 14'd121;
            {7'd11,7'd12}:		p = 14'd132;
            {7'd11,7'd13}:		p = 14'd143;
            {7'd11,7'd14}:		p = 14'd154;
            {7'd11,7'd15}:		p = 14'd165;
            {7'd11,7'd16}:		p = 14'd176;
            {7'd11,7'd17}:		p = 14'd187;
            {7'd11,7'd18}:		p = 14'd198;
            {7'd11,7'd19}:		p = 14'd209;
            {7'd11,7'd20}:		p = 14'd220;
            {7'd11,7'd21}:		p = 14'd231;
            {7'd11,7'd22}:		p = 14'd242;
            {7'd11,7'd23}:		p = 14'd253;
            {7'd11,7'd24}:		p = 14'd264;
            {7'd11,7'd25}:		p = 14'd275;
            {7'd11,7'd26}:		p = 14'd286;
            {7'd11,7'd27}:		p = 14'd297;
            {7'd11,7'd28}:		p = 14'd308;
            {7'd11,7'd29}:		p = 14'd319;
            {7'd11,7'd30}:		p = 14'd330;
            {7'd11,7'd31}:		p = 14'd341;
            {7'd11,7'd32}:		p = 14'd352;
            {7'd11,7'd33}:		p = 14'd363;
            {7'd11,7'd34}:		p = 14'd374;
            {7'd11,7'd35}:		p = 14'd385;
            {7'd11,7'd36}:		p = 14'd396;
            {7'd11,7'd37}:		p = 14'd407;
            {7'd11,7'd38}:		p = 14'd418;
            {7'd11,7'd39}:		p = 14'd429;
            {7'd11,7'd40}:		p = 14'd440;
            {7'd11,7'd41}:		p = 14'd451;
            {7'd11,7'd42}:		p = 14'd462;
            {7'd11,7'd43}:		p = 14'd473;
            {7'd11,7'd44}:		p = 14'd484;
            {7'd11,7'd45}:		p = 14'd495;
            {7'd11,7'd46}:		p = 14'd506;
            {7'd11,7'd47}:		p = 14'd517;
            {7'd11,7'd48}:		p = 14'd528;
            {7'd11,7'd49}:		p = 14'd539;
            {7'd11,7'd50}:		p = 14'd550;
            {7'd11,7'd51}:		p = 14'd561;
            {7'd11,7'd52}:		p = 14'd572;
            {7'd11,7'd53}:		p = 14'd583;
            {7'd11,7'd54}:		p = 14'd594;
            {7'd11,7'd55}:		p = 14'd605;
            {7'd11,7'd56}:		p = 14'd616;
            {7'd11,7'd57}:		p = 14'd627;
            {7'd11,7'd58}:		p = 14'd638;
            {7'd11,7'd59}:		p = 14'd649;
            {7'd11,7'd60}:		p = 14'd660;
            {7'd11,7'd61}:		p = 14'd671;
            {7'd11,7'd62}:		p = 14'd682;
            {7'd11,7'd63}:		p = 14'd693;
            {7'd11,7'd64}:		p = 14'd704;
            {7'd11,7'd65}:		p = 14'd715;
            {7'd11,7'd66}:		p = 14'd726;
            {7'd11,7'd67}:		p = 14'd737;
            {7'd11,7'd68}:		p = 14'd748;
            {7'd11,7'd69}:		p = 14'd759;
            {7'd11,7'd70}:		p = 14'd770;
            {7'd11,7'd71}:		p = 14'd781;
            {7'd11,7'd72}:		p = 14'd792;
            {7'd11,7'd73}:		p = 14'd803;
            {7'd11,7'd74}:		p = 14'd814;
            {7'd11,7'd75}:		p = 14'd825;
            {7'd11,7'd76}:		p = 14'd836;
            {7'd11,7'd77}:		p = 14'd847;
            {7'd11,7'd78}:		p = 14'd858;
            {7'd11,7'd79}:		p = 14'd869;
            {7'd11,7'd80}:		p = 14'd880;
            {7'd11,7'd81}:		p = 14'd891;
            {7'd11,7'd82}:		p = 14'd902;
            {7'd11,7'd83}:		p = 14'd913;
            {7'd11,7'd84}:		p = 14'd924;
            {7'd11,7'd85}:		p = 14'd935;
            {7'd11,7'd86}:		p = 14'd946;
            {7'd11,7'd87}:		p = 14'd957;
            {7'd11,7'd88}:		p = 14'd968;
            {7'd11,7'd89}:		p = 14'd979;
            {7'd11,7'd90}:		p = 14'd990;
            {7'd11,7'd91}:		p = 14'd1001;
            {7'd11,7'd92}:		p = 14'd1012;
            {7'd11,7'd93}:		p = 14'd1023;
            {7'd11,7'd94}:		p = 14'd1034;
            {7'd11,7'd95}:		p = 14'd1045;
            {7'd11,7'd96}:		p = 14'd1056;
            {7'd11,7'd97}:		p = 14'd1067;
            {7'd11,7'd98}:		p = 14'd1078;
            {7'd11,7'd99}:		p = 14'd1089;
            {7'd11,7'd100}:		p = 14'd1100;
            {7'd11,7'd101}:		p = 14'd1111;
            {7'd11,7'd102}:		p = 14'd1122;
            {7'd11,7'd103}:		p = 14'd1133;
            {7'd11,7'd104}:		p = 14'd1144;
            {7'd11,7'd105}:		p = 14'd1155;
            {7'd11,7'd106}:		p = 14'd1166;
            {7'd11,7'd107}:		p = 14'd1177;
            {7'd11,7'd108}:		p = 14'd1188;
            {7'd11,7'd109}:		p = 14'd1199;
            {7'd11,7'd110}:		p = 14'd1210;
            {7'd11,7'd111}:		p = 14'd1221;
            {7'd11,7'd112}:		p = 14'd1232;
            {7'd11,7'd113}:		p = 14'd1243;
            {7'd11,7'd114}:		p = 14'd1254;
            {7'd11,7'd115}:		p = 14'd1265;
            {7'd11,7'd116}:		p = 14'd1276;
            {7'd11,7'd117}:		p = 14'd1287;
            {7'd11,7'd118}:		p = 14'd1298;
            {7'd11,7'd119}:		p = 14'd1309;
            {7'd11,7'd120}:		p = 14'd1320;
            {7'd11,7'd121}:		p = 14'd1331;
            {7'd11,7'd122}:		p = 14'd1342;
            {7'd11,7'd123}:		p = 14'd1353;
            {7'd11,7'd124}:		p = 14'd1364;
            {7'd11,7'd125}:		p = 14'd1375;
            {7'd11,7'd126}:		p = 14'd1386;
            {7'd11,7'd127}:		p = 14'd1397;
            {7'd12,7'd0}:		p = 14'd0;
            {7'd12,7'd1}:		p = 14'd12;
            {7'd12,7'd2}:		p = 14'd24;
            {7'd12,7'd3}:		p = 14'd36;
            {7'd12,7'd4}:		p = 14'd48;
            {7'd12,7'd5}:		p = 14'd60;
            {7'd12,7'd6}:		p = 14'd72;
            {7'd12,7'd7}:		p = 14'd84;
            {7'd12,7'd8}:		p = 14'd96;
            {7'd12,7'd9}:		p = 14'd108;
            {7'd12,7'd10}:		p = 14'd120;
            {7'd12,7'd11}:		p = 14'd132;
            {7'd12,7'd12}:		p = 14'd144;
            {7'd12,7'd13}:		p = 14'd156;
            {7'd12,7'd14}:		p = 14'd168;
            {7'd12,7'd15}:		p = 14'd180;
            {7'd12,7'd16}:		p = 14'd192;
            {7'd12,7'd17}:		p = 14'd204;
            {7'd12,7'd18}:		p = 14'd216;
            {7'd12,7'd19}:		p = 14'd228;
            {7'd12,7'd20}:		p = 14'd240;
            {7'd12,7'd21}:		p = 14'd252;
            {7'd12,7'd22}:		p = 14'd264;
            {7'd12,7'd23}:		p = 14'd276;
            {7'd12,7'd24}:		p = 14'd288;
            {7'd12,7'd25}:		p = 14'd300;
            {7'd12,7'd26}:		p = 14'd312;
            {7'd12,7'd27}:		p = 14'd324;
            {7'd12,7'd28}:		p = 14'd336;
            {7'd12,7'd29}:		p = 14'd348;
            {7'd12,7'd30}:		p = 14'd360;
            {7'd12,7'd31}:		p = 14'd372;
            {7'd12,7'd32}:		p = 14'd384;
            {7'd12,7'd33}:		p = 14'd396;
            {7'd12,7'd34}:		p = 14'd408;
            {7'd12,7'd35}:		p = 14'd420;
            {7'd12,7'd36}:		p = 14'd432;
            {7'd12,7'd37}:		p = 14'd444;
            {7'd12,7'd38}:		p = 14'd456;
            {7'd12,7'd39}:		p = 14'd468;
            {7'd12,7'd40}:		p = 14'd480;
            {7'd12,7'd41}:		p = 14'd492;
            {7'd12,7'd42}:		p = 14'd504;
            {7'd12,7'd43}:		p = 14'd516;
            {7'd12,7'd44}:		p = 14'd528;
            {7'd12,7'd45}:		p = 14'd540;
            {7'd12,7'd46}:		p = 14'd552;
            {7'd12,7'd47}:		p = 14'd564;
            {7'd12,7'd48}:		p = 14'd576;
            {7'd12,7'd49}:		p = 14'd588;
            {7'd12,7'd50}:		p = 14'd600;
            {7'd12,7'd51}:		p = 14'd612;
            {7'd12,7'd52}:		p = 14'd624;
            {7'd12,7'd53}:		p = 14'd636;
            {7'd12,7'd54}:		p = 14'd648;
            {7'd12,7'd55}:		p = 14'd660;
            {7'd12,7'd56}:		p = 14'd672;
            {7'd12,7'd57}:		p = 14'd684;
            {7'd12,7'd58}:		p = 14'd696;
            {7'd12,7'd59}:		p = 14'd708;
            {7'd12,7'd60}:		p = 14'd720;
            {7'd12,7'd61}:		p = 14'd732;
            {7'd12,7'd62}:		p = 14'd744;
            {7'd12,7'd63}:		p = 14'd756;
            {7'd12,7'd64}:		p = 14'd768;
            {7'd12,7'd65}:		p = 14'd780;
            {7'd12,7'd66}:		p = 14'd792;
            {7'd12,7'd67}:		p = 14'd804;
            {7'd12,7'd68}:		p = 14'd816;
            {7'd12,7'd69}:		p = 14'd828;
            {7'd12,7'd70}:		p = 14'd840;
            {7'd12,7'd71}:		p = 14'd852;
            {7'd12,7'd72}:		p = 14'd864;
            {7'd12,7'd73}:		p = 14'd876;
            {7'd12,7'd74}:		p = 14'd888;
            {7'd12,7'd75}:		p = 14'd900;
            {7'd12,7'd76}:		p = 14'd912;
            {7'd12,7'd77}:		p = 14'd924;
            {7'd12,7'd78}:		p = 14'd936;
            {7'd12,7'd79}:		p = 14'd948;
            {7'd12,7'd80}:		p = 14'd960;
            {7'd12,7'd81}:		p = 14'd972;
            {7'd12,7'd82}:		p = 14'd984;
            {7'd12,7'd83}:		p = 14'd996;
            {7'd12,7'd84}:		p = 14'd1008;
            {7'd12,7'd85}:		p = 14'd1020;
            {7'd12,7'd86}:		p = 14'd1032;
            {7'd12,7'd87}:		p = 14'd1044;
            {7'd12,7'd88}:		p = 14'd1056;
            {7'd12,7'd89}:		p = 14'd1068;
            {7'd12,7'd90}:		p = 14'd1080;
            {7'd12,7'd91}:		p = 14'd1092;
            {7'd12,7'd92}:		p = 14'd1104;
            {7'd12,7'd93}:		p = 14'd1116;
            {7'd12,7'd94}:		p = 14'd1128;
            {7'd12,7'd95}:		p = 14'd1140;
            {7'd12,7'd96}:		p = 14'd1152;
            {7'd12,7'd97}:		p = 14'd1164;
            {7'd12,7'd98}:		p = 14'd1176;
            {7'd12,7'd99}:		p = 14'd1188;
            {7'd12,7'd100}:		p = 14'd1200;
            {7'd12,7'd101}:		p = 14'd1212;
            {7'd12,7'd102}:		p = 14'd1224;
            {7'd12,7'd103}:		p = 14'd1236;
            {7'd12,7'd104}:		p = 14'd1248;
            {7'd12,7'd105}:		p = 14'd1260;
            {7'd12,7'd106}:		p = 14'd1272;
            {7'd12,7'd107}:		p = 14'd1284;
            {7'd12,7'd108}:		p = 14'd1296;
            {7'd12,7'd109}:		p = 14'd1308;
            {7'd12,7'd110}:		p = 14'd1320;
            {7'd12,7'd111}:		p = 14'd1332;
            {7'd12,7'd112}:		p = 14'd1344;
            {7'd12,7'd113}:		p = 14'd1356;
            {7'd12,7'd114}:		p = 14'd1368;
            {7'd12,7'd115}:		p = 14'd1380;
            {7'd12,7'd116}:		p = 14'd1392;
            {7'd12,7'd117}:		p = 14'd1404;
            {7'd12,7'd118}:		p = 14'd1416;
            {7'd12,7'd119}:		p = 14'd1428;
            {7'd12,7'd120}:		p = 14'd1440;
            {7'd12,7'd121}:		p = 14'd1452;
            {7'd12,7'd122}:		p = 14'd1464;
            {7'd12,7'd123}:		p = 14'd1476;
            {7'd12,7'd124}:		p = 14'd1488;
            {7'd12,7'd125}:		p = 14'd1500;
            {7'd12,7'd126}:		p = 14'd1512;
            {7'd12,7'd127}:		p = 14'd1524;
            {7'd13,7'd0}:		p = 14'd0;
            {7'd13,7'd1}:		p = 14'd13;
            {7'd13,7'd2}:		p = 14'd26;
            {7'd13,7'd3}:		p = 14'd39;
            {7'd13,7'd4}:		p = 14'd52;
            {7'd13,7'd5}:		p = 14'd65;
            {7'd13,7'd6}:		p = 14'd78;
            {7'd13,7'd7}:		p = 14'd91;
            {7'd13,7'd8}:		p = 14'd104;
            {7'd13,7'd9}:		p = 14'd117;
            {7'd13,7'd10}:		p = 14'd130;
            {7'd13,7'd11}:		p = 14'd143;
            {7'd13,7'd12}:		p = 14'd156;
            {7'd13,7'd13}:		p = 14'd169;
            {7'd13,7'd14}:		p = 14'd182;
            {7'd13,7'd15}:		p = 14'd195;
            {7'd13,7'd16}:		p = 14'd208;
            {7'd13,7'd17}:		p = 14'd221;
            {7'd13,7'd18}:		p = 14'd234;
            {7'd13,7'd19}:		p = 14'd247;
            {7'd13,7'd20}:		p = 14'd260;
            {7'd13,7'd21}:		p = 14'd273;
            {7'd13,7'd22}:		p = 14'd286;
            {7'd13,7'd23}:		p = 14'd299;
            {7'd13,7'd24}:		p = 14'd312;
            {7'd13,7'd25}:		p = 14'd325;
            {7'd13,7'd26}:		p = 14'd338;
            {7'd13,7'd27}:		p = 14'd351;
            {7'd13,7'd28}:		p = 14'd364;
            {7'd13,7'd29}:		p = 14'd377;
            {7'd13,7'd30}:		p = 14'd390;
            {7'd13,7'd31}:		p = 14'd403;
            {7'd13,7'd32}:		p = 14'd416;
            {7'd13,7'd33}:		p = 14'd429;
            {7'd13,7'd34}:		p = 14'd442;
            {7'd13,7'd35}:		p = 14'd455;
            {7'd13,7'd36}:		p = 14'd468;
            {7'd13,7'd37}:		p = 14'd481;
            {7'd13,7'd38}:		p = 14'd494;
            {7'd13,7'd39}:		p = 14'd507;
            {7'd13,7'd40}:		p = 14'd520;
            {7'd13,7'd41}:		p = 14'd533;
            {7'd13,7'd42}:		p = 14'd546;
            {7'd13,7'd43}:		p = 14'd559;
            {7'd13,7'd44}:		p = 14'd572;
            {7'd13,7'd45}:		p = 14'd585;
            {7'd13,7'd46}:		p = 14'd598;
            {7'd13,7'd47}:		p = 14'd611;
            {7'd13,7'd48}:		p = 14'd624;
            {7'd13,7'd49}:		p = 14'd637;
            {7'd13,7'd50}:		p = 14'd650;
            {7'd13,7'd51}:		p = 14'd663;
            {7'd13,7'd52}:		p = 14'd676;
            {7'd13,7'd53}:		p = 14'd689;
            {7'd13,7'd54}:		p = 14'd702;
            {7'd13,7'd55}:		p = 14'd715;
            {7'd13,7'd56}:		p = 14'd728;
            {7'd13,7'd57}:		p = 14'd741;
            {7'd13,7'd58}:		p = 14'd754;
            {7'd13,7'd59}:		p = 14'd767;
            {7'd13,7'd60}:		p = 14'd780;
            {7'd13,7'd61}:		p = 14'd793;
            {7'd13,7'd62}:		p = 14'd806;
            {7'd13,7'd63}:		p = 14'd819;
            {7'd13,7'd64}:		p = 14'd832;
            {7'd13,7'd65}:		p = 14'd845;
            {7'd13,7'd66}:		p = 14'd858;
            {7'd13,7'd67}:		p = 14'd871;
            {7'd13,7'd68}:		p = 14'd884;
            {7'd13,7'd69}:		p = 14'd897;
            {7'd13,7'd70}:		p = 14'd910;
            {7'd13,7'd71}:		p = 14'd923;
            {7'd13,7'd72}:		p = 14'd936;
            {7'd13,7'd73}:		p = 14'd949;
            {7'd13,7'd74}:		p = 14'd962;
            {7'd13,7'd75}:		p = 14'd975;
            {7'd13,7'd76}:		p = 14'd988;
            {7'd13,7'd77}:		p = 14'd1001;
            {7'd13,7'd78}:		p = 14'd1014;
            {7'd13,7'd79}:		p = 14'd1027;
            {7'd13,7'd80}:		p = 14'd1040;
            {7'd13,7'd81}:		p = 14'd1053;
            {7'd13,7'd82}:		p = 14'd1066;
            {7'd13,7'd83}:		p = 14'd1079;
            {7'd13,7'd84}:		p = 14'd1092;
            {7'd13,7'd85}:		p = 14'd1105;
            {7'd13,7'd86}:		p = 14'd1118;
            {7'd13,7'd87}:		p = 14'd1131;
            {7'd13,7'd88}:		p = 14'd1144;
            {7'd13,7'd89}:		p = 14'd1157;
            {7'd13,7'd90}:		p = 14'd1170;
            {7'd13,7'd91}:		p = 14'd1183;
            {7'd13,7'd92}:		p = 14'd1196;
            {7'd13,7'd93}:		p = 14'd1209;
            {7'd13,7'd94}:		p = 14'd1222;
            {7'd13,7'd95}:		p = 14'd1235;
            {7'd13,7'd96}:		p = 14'd1248;
            {7'd13,7'd97}:		p = 14'd1261;
            {7'd13,7'd98}:		p = 14'd1274;
            {7'd13,7'd99}:		p = 14'd1287;
            {7'd13,7'd100}:		p = 14'd1300;
            {7'd13,7'd101}:		p = 14'd1313;
            {7'd13,7'd102}:		p = 14'd1326;
            {7'd13,7'd103}:		p = 14'd1339;
            {7'd13,7'd104}:		p = 14'd1352;
            {7'd13,7'd105}:		p = 14'd1365;
            {7'd13,7'd106}:		p = 14'd1378;
            {7'd13,7'd107}:		p = 14'd1391;
            {7'd13,7'd108}:		p = 14'd1404;
            {7'd13,7'd109}:		p = 14'd1417;
            {7'd13,7'd110}:		p = 14'd1430;
            {7'd13,7'd111}:		p = 14'd1443;
            {7'd13,7'd112}:		p = 14'd1456;
            {7'd13,7'd113}:		p = 14'd1469;
            {7'd13,7'd114}:		p = 14'd1482;
            {7'd13,7'd115}:		p = 14'd1495;
            {7'd13,7'd116}:		p = 14'd1508;
            {7'd13,7'd117}:		p = 14'd1521;
            {7'd13,7'd118}:		p = 14'd1534;
            {7'd13,7'd119}:		p = 14'd1547;
            {7'd13,7'd120}:		p = 14'd1560;
            {7'd13,7'd121}:		p = 14'd1573;
            {7'd13,7'd122}:		p = 14'd1586;
            {7'd13,7'd123}:		p = 14'd1599;
            {7'd13,7'd124}:		p = 14'd1612;
            {7'd13,7'd125}:		p = 14'd1625;
            {7'd13,7'd126}:		p = 14'd1638;
            {7'd13,7'd127}:		p = 14'd1651;
            {7'd14,7'd0}:		p = 14'd0;
            {7'd14,7'd1}:		p = 14'd14;
            {7'd14,7'd2}:		p = 14'd28;
            {7'd14,7'd3}:		p = 14'd42;
            {7'd14,7'd4}:		p = 14'd56;
            {7'd14,7'd5}:		p = 14'd70;
            {7'd14,7'd6}:		p = 14'd84;
            {7'd14,7'd7}:		p = 14'd98;
            {7'd14,7'd8}:		p = 14'd112;
            {7'd14,7'd9}:		p = 14'd126;
            {7'd14,7'd10}:		p = 14'd140;
            {7'd14,7'd11}:		p = 14'd154;
            {7'd14,7'd12}:		p = 14'd168;
            {7'd14,7'd13}:		p = 14'd182;
            {7'd14,7'd14}:		p = 14'd196;
            {7'd14,7'd15}:		p = 14'd210;
            {7'd14,7'd16}:		p = 14'd224;
            {7'd14,7'd17}:		p = 14'd238;
            {7'd14,7'd18}:		p = 14'd252;
            {7'd14,7'd19}:		p = 14'd266;
            {7'd14,7'd20}:		p = 14'd280;
            {7'd14,7'd21}:		p = 14'd294;
            {7'd14,7'd22}:		p = 14'd308;
            {7'd14,7'd23}:		p = 14'd322;
            {7'd14,7'd24}:		p = 14'd336;
            {7'd14,7'd25}:		p = 14'd350;
            {7'd14,7'd26}:		p = 14'd364;
            {7'd14,7'd27}:		p = 14'd378;
            {7'd14,7'd28}:		p = 14'd392;
            {7'd14,7'd29}:		p = 14'd406;
            {7'd14,7'd30}:		p = 14'd420;
            {7'd14,7'd31}:		p = 14'd434;
            {7'd14,7'd32}:		p = 14'd448;
            {7'd14,7'd33}:		p = 14'd462;
            {7'd14,7'd34}:		p = 14'd476;
            {7'd14,7'd35}:		p = 14'd490;
            {7'd14,7'd36}:		p = 14'd504;
            {7'd14,7'd37}:		p = 14'd518;
            {7'd14,7'd38}:		p = 14'd532;
            {7'd14,7'd39}:		p = 14'd546;
            {7'd14,7'd40}:		p = 14'd560;
            {7'd14,7'd41}:		p = 14'd574;
            {7'd14,7'd42}:		p = 14'd588;
            {7'd14,7'd43}:		p = 14'd602;
            {7'd14,7'd44}:		p = 14'd616;
            {7'd14,7'd45}:		p = 14'd630;
            {7'd14,7'd46}:		p = 14'd644;
            {7'd14,7'd47}:		p = 14'd658;
            {7'd14,7'd48}:		p = 14'd672;
            {7'd14,7'd49}:		p = 14'd686;
            {7'd14,7'd50}:		p = 14'd700;
            {7'd14,7'd51}:		p = 14'd714;
            {7'd14,7'd52}:		p = 14'd728;
            {7'd14,7'd53}:		p = 14'd742;
            {7'd14,7'd54}:		p = 14'd756;
            {7'd14,7'd55}:		p = 14'd770;
            {7'd14,7'd56}:		p = 14'd784;
            {7'd14,7'd57}:		p = 14'd798;
            {7'd14,7'd58}:		p = 14'd812;
            {7'd14,7'd59}:		p = 14'd826;
            {7'd14,7'd60}:		p = 14'd840;
            {7'd14,7'd61}:		p = 14'd854;
            {7'd14,7'd62}:		p = 14'd868;
            {7'd14,7'd63}:		p = 14'd882;
            {7'd14,7'd64}:		p = 14'd896;
            {7'd14,7'd65}:		p = 14'd910;
            {7'd14,7'd66}:		p = 14'd924;
            {7'd14,7'd67}:		p = 14'd938;
            {7'd14,7'd68}:		p = 14'd952;
            {7'd14,7'd69}:		p = 14'd966;
            {7'd14,7'd70}:		p = 14'd980;
            {7'd14,7'd71}:		p = 14'd994;
            {7'd14,7'd72}:		p = 14'd1008;
            {7'd14,7'd73}:		p = 14'd1022;
            {7'd14,7'd74}:		p = 14'd1036;
            {7'd14,7'd75}:		p = 14'd1050;
            {7'd14,7'd76}:		p = 14'd1064;
            {7'd14,7'd77}:		p = 14'd1078;
            {7'd14,7'd78}:		p = 14'd1092;
            {7'd14,7'd79}:		p = 14'd1106;
            {7'd14,7'd80}:		p = 14'd1120;
            {7'd14,7'd81}:		p = 14'd1134;
            {7'd14,7'd82}:		p = 14'd1148;
            {7'd14,7'd83}:		p = 14'd1162;
            {7'd14,7'd84}:		p = 14'd1176;
            {7'd14,7'd85}:		p = 14'd1190;
            {7'd14,7'd86}:		p = 14'd1204;
            {7'd14,7'd87}:		p = 14'd1218;
            {7'd14,7'd88}:		p = 14'd1232;
            {7'd14,7'd89}:		p = 14'd1246;
            {7'd14,7'd90}:		p = 14'd1260;
            {7'd14,7'd91}:		p = 14'd1274;
            {7'd14,7'd92}:		p = 14'd1288;
            {7'd14,7'd93}:		p = 14'd1302;
            {7'd14,7'd94}:		p = 14'd1316;
            {7'd14,7'd95}:		p = 14'd1330;
            {7'd14,7'd96}:		p = 14'd1344;
            {7'd14,7'd97}:		p = 14'd1358;
            {7'd14,7'd98}:		p = 14'd1372;
            {7'd14,7'd99}:		p = 14'd1386;
            {7'd14,7'd100}:		p = 14'd1400;
            {7'd14,7'd101}:		p = 14'd1414;
            {7'd14,7'd102}:		p = 14'd1428;
            {7'd14,7'd103}:		p = 14'd1442;
            {7'd14,7'd104}:		p = 14'd1456;
            {7'd14,7'd105}:		p = 14'd1470;
            {7'd14,7'd106}:		p = 14'd1484;
            {7'd14,7'd107}:		p = 14'd1498;
            {7'd14,7'd108}:		p = 14'd1512;
            {7'd14,7'd109}:		p = 14'd1526;
            {7'd14,7'd110}:		p = 14'd1540;
            {7'd14,7'd111}:		p = 14'd1554;
            {7'd14,7'd112}:		p = 14'd1568;
            {7'd14,7'd113}:		p = 14'd1582;
            {7'd14,7'd114}:		p = 14'd1596;
            {7'd14,7'd115}:		p = 14'd1610;
            {7'd14,7'd116}:		p = 14'd1624;
            {7'd14,7'd117}:		p = 14'd1638;
            {7'd14,7'd118}:		p = 14'd1652;
            {7'd14,7'd119}:		p = 14'd1666;
            {7'd14,7'd120}:		p = 14'd1680;
            {7'd14,7'd121}:		p = 14'd1694;
            {7'd14,7'd122}:		p = 14'd1708;
            {7'd14,7'd123}:		p = 14'd1722;
            {7'd14,7'd124}:		p = 14'd1736;
            {7'd14,7'd125}:		p = 14'd1750;
            {7'd14,7'd126}:		p = 14'd1764;
            {7'd14,7'd127}:		p = 14'd1778;
            {7'd15,7'd0}:		p = 14'd0;
            {7'd15,7'd1}:		p = 14'd15;
            {7'd15,7'd2}:		p = 14'd30;
            {7'd15,7'd3}:		p = 14'd45;
            {7'd15,7'd4}:		p = 14'd60;
            {7'd15,7'd5}:		p = 14'd75;
            {7'd15,7'd6}:		p = 14'd90;
            {7'd15,7'd7}:		p = 14'd105;
            {7'd15,7'd8}:		p = 14'd120;
            {7'd15,7'd9}:		p = 14'd135;
            {7'd15,7'd10}:		p = 14'd150;
            {7'd15,7'd11}:		p = 14'd165;
            {7'd15,7'd12}:		p = 14'd180;
            {7'd15,7'd13}:		p = 14'd195;
            {7'd15,7'd14}:		p = 14'd210;
            {7'd15,7'd15}:		p = 14'd225;
            {7'd15,7'd16}:		p = 14'd240;
            {7'd15,7'd17}:		p = 14'd255;
            {7'd15,7'd18}:		p = 14'd270;
            {7'd15,7'd19}:		p = 14'd285;
            {7'd15,7'd20}:		p = 14'd300;
            {7'd15,7'd21}:		p = 14'd315;
            {7'd15,7'd22}:		p = 14'd330;
            {7'd15,7'd23}:		p = 14'd345;
            {7'd15,7'd24}:		p = 14'd360;
            {7'd15,7'd25}:		p = 14'd375;
            {7'd15,7'd26}:		p = 14'd390;
            {7'd15,7'd27}:		p = 14'd405;
            {7'd15,7'd28}:		p = 14'd420;
            {7'd15,7'd29}:		p = 14'd435;
            {7'd15,7'd30}:		p = 14'd450;
            {7'd15,7'd31}:		p = 14'd465;
            {7'd15,7'd32}:		p = 14'd480;
            {7'd15,7'd33}:		p = 14'd495;
            {7'd15,7'd34}:		p = 14'd510;
            {7'd15,7'd35}:		p = 14'd525;
            {7'd15,7'd36}:		p = 14'd540;
            {7'd15,7'd37}:		p = 14'd555;
            {7'd15,7'd38}:		p = 14'd570;
            {7'd15,7'd39}:		p = 14'd585;
            {7'd15,7'd40}:		p = 14'd600;
            {7'd15,7'd41}:		p = 14'd615;
            {7'd15,7'd42}:		p = 14'd630;
            {7'd15,7'd43}:		p = 14'd645;
            {7'd15,7'd44}:		p = 14'd660;
            {7'd15,7'd45}:		p = 14'd675;
            {7'd15,7'd46}:		p = 14'd690;
            {7'd15,7'd47}:		p = 14'd705;
            {7'd15,7'd48}:		p = 14'd720;
            {7'd15,7'd49}:		p = 14'd735;
            {7'd15,7'd50}:		p = 14'd750;
            {7'd15,7'd51}:		p = 14'd765;
            {7'd15,7'd52}:		p = 14'd780;
            {7'd15,7'd53}:		p = 14'd795;
            {7'd15,7'd54}:		p = 14'd810;
            {7'd15,7'd55}:		p = 14'd825;
            {7'd15,7'd56}:		p = 14'd840;
            {7'd15,7'd57}:		p = 14'd855;
            {7'd15,7'd58}:		p = 14'd870;
            {7'd15,7'd59}:		p = 14'd885;
            {7'd15,7'd60}:		p = 14'd900;
            {7'd15,7'd61}:		p = 14'd915;
            {7'd15,7'd62}:		p = 14'd930;
            {7'd15,7'd63}:		p = 14'd945;
            {7'd15,7'd64}:		p = 14'd960;
            {7'd15,7'd65}:		p = 14'd975;
            {7'd15,7'd66}:		p = 14'd990;
            {7'd15,7'd67}:		p = 14'd1005;
            {7'd15,7'd68}:		p = 14'd1020;
            {7'd15,7'd69}:		p = 14'd1035;
            {7'd15,7'd70}:		p = 14'd1050;
            {7'd15,7'd71}:		p = 14'd1065;
            {7'd15,7'd72}:		p = 14'd1080;
            {7'd15,7'd73}:		p = 14'd1095;
            {7'd15,7'd74}:		p = 14'd1110;
            {7'd15,7'd75}:		p = 14'd1125;
            {7'd15,7'd76}:		p = 14'd1140;
            {7'd15,7'd77}:		p = 14'd1155;
            {7'd15,7'd78}:		p = 14'd1170;
            {7'd15,7'd79}:		p = 14'd1185;
            {7'd15,7'd80}:		p = 14'd1200;
            {7'd15,7'd81}:		p = 14'd1215;
            {7'd15,7'd82}:		p = 14'd1230;
            {7'd15,7'd83}:		p = 14'd1245;
            {7'd15,7'd84}:		p = 14'd1260;
            {7'd15,7'd85}:		p = 14'd1275;
            {7'd15,7'd86}:		p = 14'd1290;
            {7'd15,7'd87}:		p = 14'd1305;
            {7'd15,7'd88}:		p = 14'd1320;
            {7'd15,7'd89}:		p = 14'd1335;
            {7'd15,7'd90}:		p = 14'd1350;
            {7'd15,7'd91}:		p = 14'd1365;
            {7'd15,7'd92}:		p = 14'd1380;
            {7'd15,7'd93}:		p = 14'd1395;
            {7'd15,7'd94}:		p = 14'd1410;
            {7'd15,7'd95}:		p = 14'd1425;
            {7'd15,7'd96}:		p = 14'd1440;
            {7'd15,7'd97}:		p = 14'd1455;
            {7'd15,7'd98}:		p = 14'd1470;
            {7'd15,7'd99}:		p = 14'd1485;
            {7'd15,7'd100}:		p = 14'd1500;
            {7'd15,7'd101}:		p = 14'd1515;
            {7'd15,7'd102}:		p = 14'd1530;
            {7'd15,7'd103}:		p = 14'd1545;
            {7'd15,7'd104}:		p = 14'd1560;
            {7'd15,7'd105}:		p = 14'd1575;
            {7'd15,7'd106}:		p = 14'd1590;
            {7'd15,7'd107}:		p = 14'd1605;
            {7'd15,7'd108}:		p = 14'd1620;
            {7'd15,7'd109}:		p = 14'd1635;
            {7'd15,7'd110}:		p = 14'd1650;
            {7'd15,7'd111}:		p = 14'd1665;
            {7'd15,7'd112}:		p = 14'd1680;
            {7'd15,7'd113}:		p = 14'd1695;
            {7'd15,7'd114}:		p = 14'd1710;
            {7'd15,7'd115}:		p = 14'd1725;
            {7'd15,7'd116}:		p = 14'd1740;
            {7'd15,7'd117}:		p = 14'd1755;
            {7'd15,7'd118}:		p = 14'd1770;
            {7'd15,7'd119}:		p = 14'd1785;
            {7'd15,7'd120}:		p = 14'd1800;
            {7'd15,7'd121}:		p = 14'd1815;
            {7'd15,7'd122}:		p = 14'd1830;
            {7'd15,7'd123}:		p = 14'd1845;
            {7'd15,7'd124}:		p = 14'd1860;
            {7'd15,7'd125}:		p = 14'd1875;
            {7'd15,7'd126}:		p = 14'd1890;
            {7'd15,7'd127}:		p = 14'd1905;
            {7'd16,7'd0}:		p = 14'd0;
            {7'd16,7'd1}:		p = 14'd16;
            {7'd16,7'd2}:		p = 14'd32;
            {7'd16,7'd3}:		p = 14'd48;
            {7'd16,7'd4}:		p = 14'd64;
            {7'd16,7'd5}:		p = 14'd80;
            {7'd16,7'd6}:		p = 14'd96;
            {7'd16,7'd7}:		p = 14'd112;
            {7'd16,7'd8}:		p = 14'd128;
            {7'd16,7'd9}:		p = 14'd144;
            {7'd16,7'd10}:		p = 14'd160;
            {7'd16,7'd11}:		p = 14'd176;
            {7'd16,7'd12}:		p = 14'd192;
            {7'd16,7'd13}:		p = 14'd208;
            {7'd16,7'd14}:		p = 14'd224;
            {7'd16,7'd15}:		p = 14'd240;
            {7'd16,7'd16}:		p = 14'd256;
            {7'd16,7'd17}:		p = 14'd272;
            {7'd16,7'd18}:		p = 14'd288;
            {7'd16,7'd19}:		p = 14'd304;
            {7'd16,7'd20}:		p = 14'd320;
            {7'd16,7'd21}:		p = 14'd336;
            {7'd16,7'd22}:		p = 14'd352;
            {7'd16,7'd23}:		p = 14'd368;
            {7'd16,7'd24}:		p = 14'd384;
            {7'd16,7'd25}:		p = 14'd400;
            {7'd16,7'd26}:		p = 14'd416;
            {7'd16,7'd27}:		p = 14'd432;
            {7'd16,7'd28}:		p = 14'd448;
            {7'd16,7'd29}:		p = 14'd464;
            {7'd16,7'd30}:		p = 14'd480;
            {7'd16,7'd31}:		p = 14'd496;
            {7'd16,7'd32}:		p = 14'd512;
            {7'd16,7'd33}:		p = 14'd528;
            {7'd16,7'd34}:		p = 14'd544;
            {7'd16,7'd35}:		p = 14'd560;
            {7'd16,7'd36}:		p = 14'd576;
            {7'd16,7'd37}:		p = 14'd592;
            {7'd16,7'd38}:		p = 14'd608;
            {7'd16,7'd39}:		p = 14'd624;
            {7'd16,7'd40}:		p = 14'd640;
            {7'd16,7'd41}:		p = 14'd656;
            {7'd16,7'd42}:		p = 14'd672;
            {7'd16,7'd43}:		p = 14'd688;
            {7'd16,7'd44}:		p = 14'd704;
            {7'd16,7'd45}:		p = 14'd720;
            {7'd16,7'd46}:		p = 14'd736;
            {7'd16,7'd47}:		p = 14'd752;
            {7'd16,7'd48}:		p = 14'd768;
            {7'd16,7'd49}:		p = 14'd784;
            {7'd16,7'd50}:		p = 14'd800;
            {7'd16,7'd51}:		p = 14'd816;
            {7'd16,7'd52}:		p = 14'd832;
            {7'd16,7'd53}:		p = 14'd848;
            {7'd16,7'd54}:		p = 14'd864;
            {7'd16,7'd55}:		p = 14'd880;
            {7'd16,7'd56}:		p = 14'd896;
            {7'd16,7'd57}:		p = 14'd912;
            {7'd16,7'd58}:		p = 14'd928;
            {7'd16,7'd59}:		p = 14'd944;
            {7'd16,7'd60}:		p = 14'd960;
            {7'd16,7'd61}:		p = 14'd976;
            {7'd16,7'd62}:		p = 14'd992;
            {7'd16,7'd63}:		p = 14'd1008;
            {7'd16,7'd64}:		p = 14'd1024;
            {7'd16,7'd65}:		p = 14'd1040;
            {7'd16,7'd66}:		p = 14'd1056;
            {7'd16,7'd67}:		p = 14'd1072;
            {7'd16,7'd68}:		p = 14'd1088;
            {7'd16,7'd69}:		p = 14'd1104;
            {7'd16,7'd70}:		p = 14'd1120;
            {7'd16,7'd71}:		p = 14'd1136;
            {7'd16,7'd72}:		p = 14'd1152;
            {7'd16,7'd73}:		p = 14'd1168;
            {7'd16,7'd74}:		p = 14'd1184;
            {7'd16,7'd75}:		p = 14'd1200;
            {7'd16,7'd76}:		p = 14'd1216;
            {7'd16,7'd77}:		p = 14'd1232;
            {7'd16,7'd78}:		p = 14'd1248;
            {7'd16,7'd79}:		p = 14'd1264;
            {7'd16,7'd80}:		p = 14'd1280;
            {7'd16,7'd81}:		p = 14'd1296;
            {7'd16,7'd82}:		p = 14'd1312;
            {7'd16,7'd83}:		p = 14'd1328;
            {7'd16,7'd84}:		p = 14'd1344;
            {7'd16,7'd85}:		p = 14'd1360;
            {7'd16,7'd86}:		p = 14'd1376;
            {7'd16,7'd87}:		p = 14'd1392;
            {7'd16,7'd88}:		p = 14'd1408;
            {7'd16,7'd89}:		p = 14'd1424;
            {7'd16,7'd90}:		p = 14'd1440;
            {7'd16,7'd91}:		p = 14'd1456;
            {7'd16,7'd92}:		p = 14'd1472;
            {7'd16,7'd93}:		p = 14'd1488;
            {7'd16,7'd94}:		p = 14'd1504;
            {7'd16,7'd95}:		p = 14'd1520;
            {7'd16,7'd96}:		p = 14'd1536;
            {7'd16,7'd97}:		p = 14'd1552;
            {7'd16,7'd98}:		p = 14'd1568;
            {7'd16,7'd99}:		p = 14'd1584;
            {7'd16,7'd100}:		p = 14'd1600;
            {7'd16,7'd101}:		p = 14'd1616;
            {7'd16,7'd102}:		p = 14'd1632;
            {7'd16,7'd103}:		p = 14'd1648;
            {7'd16,7'd104}:		p = 14'd1664;
            {7'd16,7'd105}:		p = 14'd1680;
            {7'd16,7'd106}:		p = 14'd1696;
            {7'd16,7'd107}:		p = 14'd1712;
            {7'd16,7'd108}:		p = 14'd1728;
            {7'd16,7'd109}:		p = 14'd1744;
            {7'd16,7'd110}:		p = 14'd1760;
            {7'd16,7'd111}:		p = 14'd1776;
            {7'd16,7'd112}:		p = 14'd1792;
            {7'd16,7'd113}:		p = 14'd1808;
            {7'd16,7'd114}:		p = 14'd1824;
            {7'd16,7'd115}:		p = 14'd1840;
            {7'd16,7'd116}:		p = 14'd1856;
            {7'd16,7'd117}:		p = 14'd1872;
            {7'd16,7'd118}:		p = 14'd1888;
            {7'd16,7'd119}:		p = 14'd1904;
            {7'd16,7'd120}:		p = 14'd1920;
            {7'd16,7'd121}:		p = 14'd1936;
            {7'd16,7'd122}:		p = 14'd1952;
            {7'd16,7'd123}:		p = 14'd1968;
            {7'd16,7'd124}:		p = 14'd1984;
            {7'd16,7'd125}:		p = 14'd2000;
            {7'd16,7'd126}:		p = 14'd2016;
            {7'd16,7'd127}:		p = 14'd2032;
            {7'd17,7'd0}:		p = 14'd0;
            {7'd17,7'd1}:		p = 14'd17;
            {7'd17,7'd2}:		p = 14'd34;
            {7'd17,7'd3}:		p = 14'd51;
            {7'd17,7'd4}:		p = 14'd68;
            {7'd17,7'd5}:		p = 14'd85;
            {7'd17,7'd6}:		p = 14'd102;
            {7'd17,7'd7}:		p = 14'd119;
            {7'd17,7'd8}:		p = 14'd136;
            {7'd17,7'd9}:		p = 14'd153;
            {7'd17,7'd10}:		p = 14'd170;
            {7'd17,7'd11}:		p = 14'd187;
            {7'd17,7'd12}:		p = 14'd204;
            {7'd17,7'd13}:		p = 14'd221;
            {7'd17,7'd14}:		p = 14'd238;
            {7'd17,7'd15}:		p = 14'd255;
            {7'd17,7'd16}:		p = 14'd272;
            {7'd17,7'd17}:		p = 14'd289;
            {7'd17,7'd18}:		p = 14'd306;
            {7'd17,7'd19}:		p = 14'd323;
            {7'd17,7'd20}:		p = 14'd340;
            {7'd17,7'd21}:		p = 14'd357;
            {7'd17,7'd22}:		p = 14'd374;
            {7'd17,7'd23}:		p = 14'd391;
            {7'd17,7'd24}:		p = 14'd408;
            {7'd17,7'd25}:		p = 14'd425;
            {7'd17,7'd26}:		p = 14'd442;
            {7'd17,7'd27}:		p = 14'd459;
            {7'd17,7'd28}:		p = 14'd476;
            {7'd17,7'd29}:		p = 14'd493;
            {7'd17,7'd30}:		p = 14'd510;
            {7'd17,7'd31}:		p = 14'd527;
            {7'd17,7'd32}:		p = 14'd544;
            {7'd17,7'd33}:		p = 14'd561;
            {7'd17,7'd34}:		p = 14'd578;
            {7'd17,7'd35}:		p = 14'd595;
            {7'd17,7'd36}:		p = 14'd612;
            {7'd17,7'd37}:		p = 14'd629;
            {7'd17,7'd38}:		p = 14'd646;
            {7'd17,7'd39}:		p = 14'd663;
            {7'd17,7'd40}:		p = 14'd680;
            {7'd17,7'd41}:		p = 14'd697;
            {7'd17,7'd42}:		p = 14'd714;
            {7'd17,7'd43}:		p = 14'd731;
            {7'd17,7'd44}:		p = 14'd748;
            {7'd17,7'd45}:		p = 14'd765;
            {7'd17,7'd46}:		p = 14'd782;
            {7'd17,7'd47}:		p = 14'd799;
            {7'd17,7'd48}:		p = 14'd816;
            {7'd17,7'd49}:		p = 14'd833;
            {7'd17,7'd50}:		p = 14'd850;
            {7'd17,7'd51}:		p = 14'd867;
            {7'd17,7'd52}:		p = 14'd884;
            {7'd17,7'd53}:		p = 14'd901;
            {7'd17,7'd54}:		p = 14'd918;
            {7'd17,7'd55}:		p = 14'd935;
            {7'd17,7'd56}:		p = 14'd952;
            {7'd17,7'd57}:		p = 14'd969;
            {7'd17,7'd58}:		p = 14'd986;
            {7'd17,7'd59}:		p = 14'd1003;
            {7'd17,7'd60}:		p = 14'd1020;
            {7'd17,7'd61}:		p = 14'd1037;
            {7'd17,7'd62}:		p = 14'd1054;
            {7'd17,7'd63}:		p = 14'd1071;
            {7'd17,7'd64}:		p = 14'd1088;
            {7'd17,7'd65}:		p = 14'd1105;
            {7'd17,7'd66}:		p = 14'd1122;
            {7'd17,7'd67}:		p = 14'd1139;
            {7'd17,7'd68}:		p = 14'd1156;
            {7'd17,7'd69}:		p = 14'd1173;
            {7'd17,7'd70}:		p = 14'd1190;
            {7'd17,7'd71}:		p = 14'd1207;
            {7'd17,7'd72}:		p = 14'd1224;
            {7'd17,7'd73}:		p = 14'd1241;
            {7'd17,7'd74}:		p = 14'd1258;
            {7'd17,7'd75}:		p = 14'd1275;
            {7'd17,7'd76}:		p = 14'd1292;
            {7'd17,7'd77}:		p = 14'd1309;
            {7'd17,7'd78}:		p = 14'd1326;
            {7'd17,7'd79}:		p = 14'd1343;
            {7'd17,7'd80}:		p = 14'd1360;
            {7'd17,7'd81}:		p = 14'd1377;
            {7'd17,7'd82}:		p = 14'd1394;
            {7'd17,7'd83}:		p = 14'd1411;
            {7'd17,7'd84}:		p = 14'd1428;
            {7'd17,7'd85}:		p = 14'd1445;
            {7'd17,7'd86}:		p = 14'd1462;
            {7'd17,7'd87}:		p = 14'd1479;
            {7'd17,7'd88}:		p = 14'd1496;
            {7'd17,7'd89}:		p = 14'd1513;
            {7'd17,7'd90}:		p = 14'd1530;
            {7'd17,7'd91}:		p = 14'd1547;
            {7'd17,7'd92}:		p = 14'd1564;
            {7'd17,7'd93}:		p = 14'd1581;
            {7'd17,7'd94}:		p = 14'd1598;
            {7'd17,7'd95}:		p = 14'd1615;
            {7'd17,7'd96}:		p = 14'd1632;
            {7'd17,7'd97}:		p = 14'd1649;
            {7'd17,7'd98}:		p = 14'd1666;
            {7'd17,7'd99}:		p = 14'd1683;
            {7'd17,7'd100}:		p = 14'd1700;
            {7'd17,7'd101}:		p = 14'd1717;
            {7'd17,7'd102}:		p = 14'd1734;
            {7'd17,7'd103}:		p = 14'd1751;
            {7'd17,7'd104}:		p = 14'd1768;
            {7'd17,7'd105}:		p = 14'd1785;
            {7'd17,7'd106}:		p = 14'd1802;
            {7'd17,7'd107}:		p = 14'd1819;
            {7'd17,7'd108}:		p = 14'd1836;
            {7'd17,7'd109}:		p = 14'd1853;
            {7'd17,7'd110}:		p = 14'd1870;
            {7'd17,7'd111}:		p = 14'd1887;
            {7'd17,7'd112}:		p = 14'd1904;
            {7'd17,7'd113}:		p = 14'd1921;
            {7'd17,7'd114}:		p = 14'd1938;
            {7'd17,7'd115}:		p = 14'd1955;
            {7'd17,7'd116}:		p = 14'd1972;
            {7'd17,7'd117}:		p = 14'd1989;
            {7'd17,7'd118}:		p = 14'd2006;
            {7'd17,7'd119}:		p = 14'd2023;
            {7'd17,7'd120}:		p = 14'd2040;
            {7'd17,7'd121}:		p = 14'd2057;
            {7'd17,7'd122}:		p = 14'd2074;
            {7'd17,7'd123}:		p = 14'd2091;
            {7'd17,7'd124}:		p = 14'd2108;
            {7'd17,7'd125}:		p = 14'd2125;
            {7'd17,7'd126}:		p = 14'd2142;
            {7'd17,7'd127}:		p = 14'd2159;
            {7'd18,7'd0}:		p = 14'd0;
            {7'd18,7'd1}:		p = 14'd18;
            {7'd18,7'd2}:		p = 14'd36;
            {7'd18,7'd3}:		p = 14'd54;
            {7'd18,7'd4}:		p = 14'd72;
            {7'd18,7'd5}:		p = 14'd90;
            {7'd18,7'd6}:		p = 14'd108;
            {7'd18,7'd7}:		p = 14'd126;
            {7'd18,7'd8}:		p = 14'd144;
            {7'd18,7'd9}:		p = 14'd162;
            {7'd18,7'd10}:		p = 14'd180;
            {7'd18,7'd11}:		p = 14'd198;
            {7'd18,7'd12}:		p = 14'd216;
            {7'd18,7'd13}:		p = 14'd234;
            {7'd18,7'd14}:		p = 14'd252;
            {7'd18,7'd15}:		p = 14'd270;
            {7'd18,7'd16}:		p = 14'd288;
            {7'd18,7'd17}:		p = 14'd306;
            {7'd18,7'd18}:		p = 14'd324;
            {7'd18,7'd19}:		p = 14'd342;
            {7'd18,7'd20}:		p = 14'd360;
            {7'd18,7'd21}:		p = 14'd378;
            {7'd18,7'd22}:		p = 14'd396;
            {7'd18,7'd23}:		p = 14'd414;
            {7'd18,7'd24}:		p = 14'd432;
            {7'd18,7'd25}:		p = 14'd450;
            {7'd18,7'd26}:		p = 14'd468;
            {7'd18,7'd27}:		p = 14'd486;
            {7'd18,7'd28}:		p = 14'd504;
            {7'd18,7'd29}:		p = 14'd522;
            {7'd18,7'd30}:		p = 14'd540;
            {7'd18,7'd31}:		p = 14'd558;
            {7'd18,7'd32}:		p = 14'd576;
            {7'd18,7'd33}:		p = 14'd594;
            {7'd18,7'd34}:		p = 14'd612;
            {7'd18,7'd35}:		p = 14'd630;
            {7'd18,7'd36}:		p = 14'd648;
            {7'd18,7'd37}:		p = 14'd666;
            {7'd18,7'd38}:		p = 14'd684;
            {7'd18,7'd39}:		p = 14'd702;
            {7'd18,7'd40}:		p = 14'd720;
            {7'd18,7'd41}:		p = 14'd738;
            {7'd18,7'd42}:		p = 14'd756;
            {7'd18,7'd43}:		p = 14'd774;
            {7'd18,7'd44}:		p = 14'd792;
            {7'd18,7'd45}:		p = 14'd810;
            {7'd18,7'd46}:		p = 14'd828;
            {7'd18,7'd47}:		p = 14'd846;
            {7'd18,7'd48}:		p = 14'd864;
            {7'd18,7'd49}:		p = 14'd882;
            {7'd18,7'd50}:		p = 14'd900;
            {7'd18,7'd51}:		p = 14'd918;
            {7'd18,7'd52}:		p = 14'd936;
            {7'd18,7'd53}:		p = 14'd954;
            {7'd18,7'd54}:		p = 14'd972;
            {7'd18,7'd55}:		p = 14'd990;
            {7'd18,7'd56}:		p = 14'd1008;
            {7'd18,7'd57}:		p = 14'd1026;
            {7'd18,7'd58}:		p = 14'd1044;
            {7'd18,7'd59}:		p = 14'd1062;
            {7'd18,7'd60}:		p = 14'd1080;
            {7'd18,7'd61}:		p = 14'd1098;
            {7'd18,7'd62}:		p = 14'd1116;
            {7'd18,7'd63}:		p = 14'd1134;
            {7'd18,7'd64}:		p = 14'd1152;
            {7'd18,7'd65}:		p = 14'd1170;
            {7'd18,7'd66}:		p = 14'd1188;
            {7'd18,7'd67}:		p = 14'd1206;
            {7'd18,7'd68}:		p = 14'd1224;
            {7'd18,7'd69}:		p = 14'd1242;
            {7'd18,7'd70}:		p = 14'd1260;
            {7'd18,7'd71}:		p = 14'd1278;
            {7'd18,7'd72}:		p = 14'd1296;
            {7'd18,7'd73}:		p = 14'd1314;
            {7'd18,7'd74}:		p = 14'd1332;
            {7'd18,7'd75}:		p = 14'd1350;
            {7'd18,7'd76}:		p = 14'd1368;
            {7'd18,7'd77}:		p = 14'd1386;
            {7'd18,7'd78}:		p = 14'd1404;
            {7'd18,7'd79}:		p = 14'd1422;
            {7'd18,7'd80}:		p = 14'd1440;
            {7'd18,7'd81}:		p = 14'd1458;
            {7'd18,7'd82}:		p = 14'd1476;
            {7'd18,7'd83}:		p = 14'd1494;
            {7'd18,7'd84}:		p = 14'd1512;
            {7'd18,7'd85}:		p = 14'd1530;
            {7'd18,7'd86}:		p = 14'd1548;
            {7'd18,7'd87}:		p = 14'd1566;
            {7'd18,7'd88}:		p = 14'd1584;
            {7'd18,7'd89}:		p = 14'd1602;
            {7'd18,7'd90}:		p = 14'd1620;
            {7'd18,7'd91}:		p = 14'd1638;
            {7'd18,7'd92}:		p = 14'd1656;
            {7'd18,7'd93}:		p = 14'd1674;
            {7'd18,7'd94}:		p = 14'd1692;
            {7'd18,7'd95}:		p = 14'd1710;
            {7'd18,7'd96}:		p = 14'd1728;
            {7'd18,7'd97}:		p = 14'd1746;
            {7'd18,7'd98}:		p = 14'd1764;
            {7'd18,7'd99}:		p = 14'd1782;
            {7'd18,7'd100}:		p = 14'd1800;
            {7'd18,7'd101}:		p = 14'd1818;
            {7'd18,7'd102}:		p = 14'd1836;
            {7'd18,7'd103}:		p = 14'd1854;
            {7'd18,7'd104}:		p = 14'd1872;
            {7'd18,7'd105}:		p = 14'd1890;
            {7'd18,7'd106}:		p = 14'd1908;
            {7'd18,7'd107}:		p = 14'd1926;
            {7'd18,7'd108}:		p = 14'd1944;
            {7'd18,7'd109}:		p = 14'd1962;
            {7'd18,7'd110}:		p = 14'd1980;
            {7'd18,7'd111}:		p = 14'd1998;
            {7'd18,7'd112}:		p = 14'd2016;
            {7'd18,7'd113}:		p = 14'd2034;
            {7'd18,7'd114}:		p = 14'd2052;
            {7'd18,7'd115}:		p = 14'd2070;
            {7'd18,7'd116}:		p = 14'd2088;
            {7'd18,7'd117}:		p = 14'd2106;
            {7'd18,7'd118}:		p = 14'd2124;
            {7'd18,7'd119}:		p = 14'd2142;
            {7'd18,7'd120}:		p = 14'd2160;
            {7'd18,7'd121}:		p = 14'd2178;
            {7'd18,7'd122}:		p = 14'd2196;
            {7'd18,7'd123}:		p = 14'd2214;
            {7'd18,7'd124}:		p = 14'd2232;
            {7'd18,7'd125}:		p = 14'd2250;
            {7'd18,7'd126}:		p = 14'd2268;
            {7'd18,7'd127}:		p = 14'd2286;
            {7'd19,7'd0}:		p = 14'd0;
            {7'd19,7'd1}:		p = 14'd19;
            {7'd19,7'd2}:		p = 14'd38;
            {7'd19,7'd3}:		p = 14'd57;
            {7'd19,7'd4}:		p = 14'd76;
            {7'd19,7'd5}:		p = 14'd95;
            {7'd19,7'd6}:		p = 14'd114;
            {7'd19,7'd7}:		p = 14'd133;
            {7'd19,7'd8}:		p = 14'd152;
            {7'd19,7'd9}:		p = 14'd171;
            {7'd19,7'd10}:		p = 14'd190;
            {7'd19,7'd11}:		p = 14'd209;
            {7'd19,7'd12}:		p = 14'd228;
            {7'd19,7'd13}:		p = 14'd247;
            {7'd19,7'd14}:		p = 14'd266;
            {7'd19,7'd15}:		p = 14'd285;
            {7'd19,7'd16}:		p = 14'd304;
            {7'd19,7'd17}:		p = 14'd323;
            {7'd19,7'd18}:		p = 14'd342;
            {7'd19,7'd19}:		p = 14'd361;
            {7'd19,7'd20}:		p = 14'd380;
            {7'd19,7'd21}:		p = 14'd399;
            {7'd19,7'd22}:		p = 14'd418;
            {7'd19,7'd23}:		p = 14'd437;
            {7'd19,7'd24}:		p = 14'd456;
            {7'd19,7'd25}:		p = 14'd475;
            {7'd19,7'd26}:		p = 14'd494;
            {7'd19,7'd27}:		p = 14'd513;
            {7'd19,7'd28}:		p = 14'd532;
            {7'd19,7'd29}:		p = 14'd551;
            {7'd19,7'd30}:		p = 14'd570;
            {7'd19,7'd31}:		p = 14'd589;
            {7'd19,7'd32}:		p = 14'd608;
            {7'd19,7'd33}:		p = 14'd627;
            {7'd19,7'd34}:		p = 14'd646;
            {7'd19,7'd35}:		p = 14'd665;
            {7'd19,7'd36}:		p = 14'd684;
            {7'd19,7'd37}:		p = 14'd703;
            {7'd19,7'd38}:		p = 14'd722;
            {7'd19,7'd39}:		p = 14'd741;
            {7'd19,7'd40}:		p = 14'd760;
            {7'd19,7'd41}:		p = 14'd779;
            {7'd19,7'd42}:		p = 14'd798;
            {7'd19,7'd43}:		p = 14'd817;
            {7'd19,7'd44}:		p = 14'd836;
            {7'd19,7'd45}:		p = 14'd855;
            {7'd19,7'd46}:		p = 14'd874;
            {7'd19,7'd47}:		p = 14'd893;
            {7'd19,7'd48}:		p = 14'd912;
            {7'd19,7'd49}:		p = 14'd931;
            {7'd19,7'd50}:		p = 14'd950;
            {7'd19,7'd51}:		p = 14'd969;
            {7'd19,7'd52}:		p = 14'd988;
            {7'd19,7'd53}:		p = 14'd1007;
            {7'd19,7'd54}:		p = 14'd1026;
            {7'd19,7'd55}:		p = 14'd1045;
            {7'd19,7'd56}:		p = 14'd1064;
            {7'd19,7'd57}:		p = 14'd1083;
            {7'd19,7'd58}:		p = 14'd1102;
            {7'd19,7'd59}:		p = 14'd1121;
            {7'd19,7'd60}:		p = 14'd1140;
            {7'd19,7'd61}:		p = 14'd1159;
            {7'd19,7'd62}:		p = 14'd1178;
            {7'd19,7'd63}:		p = 14'd1197;
            {7'd19,7'd64}:		p = 14'd1216;
            {7'd19,7'd65}:		p = 14'd1235;
            {7'd19,7'd66}:		p = 14'd1254;
            {7'd19,7'd67}:		p = 14'd1273;
            {7'd19,7'd68}:		p = 14'd1292;
            {7'd19,7'd69}:		p = 14'd1311;
            {7'd19,7'd70}:		p = 14'd1330;
            {7'd19,7'd71}:		p = 14'd1349;
            {7'd19,7'd72}:		p = 14'd1368;
            {7'd19,7'd73}:		p = 14'd1387;
            {7'd19,7'd74}:		p = 14'd1406;
            {7'd19,7'd75}:		p = 14'd1425;
            {7'd19,7'd76}:		p = 14'd1444;
            {7'd19,7'd77}:		p = 14'd1463;
            {7'd19,7'd78}:		p = 14'd1482;
            {7'd19,7'd79}:		p = 14'd1501;
            {7'd19,7'd80}:		p = 14'd1520;
            {7'd19,7'd81}:		p = 14'd1539;
            {7'd19,7'd82}:		p = 14'd1558;
            {7'd19,7'd83}:		p = 14'd1577;
            {7'd19,7'd84}:		p = 14'd1596;
            {7'd19,7'd85}:		p = 14'd1615;
            {7'd19,7'd86}:		p = 14'd1634;
            {7'd19,7'd87}:		p = 14'd1653;
            {7'd19,7'd88}:		p = 14'd1672;
            {7'd19,7'd89}:		p = 14'd1691;
            {7'd19,7'd90}:		p = 14'd1710;
            {7'd19,7'd91}:		p = 14'd1729;
            {7'd19,7'd92}:		p = 14'd1748;
            {7'd19,7'd93}:		p = 14'd1767;
            {7'd19,7'd94}:		p = 14'd1786;
            {7'd19,7'd95}:		p = 14'd1805;
            {7'd19,7'd96}:		p = 14'd1824;
            {7'd19,7'd97}:		p = 14'd1843;
            {7'd19,7'd98}:		p = 14'd1862;
            {7'd19,7'd99}:		p = 14'd1881;
            {7'd19,7'd100}:		p = 14'd1900;
            {7'd19,7'd101}:		p = 14'd1919;
            {7'd19,7'd102}:		p = 14'd1938;
            {7'd19,7'd103}:		p = 14'd1957;
            {7'd19,7'd104}:		p = 14'd1976;
            {7'd19,7'd105}:		p = 14'd1995;
            {7'd19,7'd106}:		p = 14'd2014;
            {7'd19,7'd107}:		p = 14'd2033;
            {7'd19,7'd108}:		p = 14'd2052;
            {7'd19,7'd109}:		p = 14'd2071;
            {7'd19,7'd110}:		p = 14'd2090;
            {7'd19,7'd111}:		p = 14'd2109;
            {7'd19,7'd112}:		p = 14'd2128;
            {7'd19,7'd113}:		p = 14'd2147;
            {7'd19,7'd114}:		p = 14'd2166;
            {7'd19,7'd115}:		p = 14'd2185;
            {7'd19,7'd116}:		p = 14'd2204;
            {7'd19,7'd117}:		p = 14'd2223;
            {7'd19,7'd118}:		p = 14'd2242;
            {7'd19,7'd119}:		p = 14'd2261;
            {7'd19,7'd120}:		p = 14'd2280;
            {7'd19,7'd121}:		p = 14'd2299;
            {7'd19,7'd122}:		p = 14'd2318;
            {7'd19,7'd123}:		p = 14'd2337;
            {7'd19,7'd124}:		p = 14'd2356;
            {7'd19,7'd125}:		p = 14'd2375;
            {7'd19,7'd126}:		p = 14'd2394;
            {7'd19,7'd127}:		p = 14'd2413;
            {7'd20,7'd0}:		p = 14'd0;
            {7'd20,7'd1}:		p = 14'd20;
            {7'd20,7'd2}:		p = 14'd40;
            {7'd20,7'd3}:		p = 14'd60;
            {7'd20,7'd4}:		p = 14'd80;
            {7'd20,7'd5}:		p = 14'd100;
            {7'd20,7'd6}:		p = 14'd120;
            {7'd20,7'd7}:		p = 14'd140;
            {7'd20,7'd8}:		p = 14'd160;
            {7'd20,7'd9}:		p = 14'd180;
            {7'd20,7'd10}:		p = 14'd200;
            {7'd20,7'd11}:		p = 14'd220;
            {7'd20,7'd12}:		p = 14'd240;
            {7'd20,7'd13}:		p = 14'd260;
            {7'd20,7'd14}:		p = 14'd280;
            {7'd20,7'd15}:		p = 14'd300;
            {7'd20,7'd16}:		p = 14'd320;
            {7'd20,7'd17}:		p = 14'd340;
            {7'd20,7'd18}:		p = 14'd360;
            {7'd20,7'd19}:		p = 14'd380;
            {7'd20,7'd20}:		p = 14'd400;
            {7'd20,7'd21}:		p = 14'd420;
            {7'd20,7'd22}:		p = 14'd440;
            {7'd20,7'd23}:		p = 14'd460;
            {7'd20,7'd24}:		p = 14'd480;
            {7'd20,7'd25}:		p = 14'd500;
            {7'd20,7'd26}:		p = 14'd520;
            {7'd20,7'd27}:		p = 14'd540;
            {7'd20,7'd28}:		p = 14'd560;
            {7'd20,7'd29}:		p = 14'd580;
            {7'd20,7'd30}:		p = 14'd600;
            {7'd20,7'd31}:		p = 14'd620;
            {7'd20,7'd32}:		p = 14'd640;
            {7'd20,7'd33}:		p = 14'd660;
            {7'd20,7'd34}:		p = 14'd680;
            {7'd20,7'd35}:		p = 14'd700;
            {7'd20,7'd36}:		p = 14'd720;
            {7'd20,7'd37}:		p = 14'd740;
            {7'd20,7'd38}:		p = 14'd760;
            {7'd20,7'd39}:		p = 14'd780;
            {7'd20,7'd40}:		p = 14'd800;
            {7'd20,7'd41}:		p = 14'd820;
            {7'd20,7'd42}:		p = 14'd840;
            {7'd20,7'd43}:		p = 14'd860;
            {7'd20,7'd44}:		p = 14'd880;
            {7'd20,7'd45}:		p = 14'd900;
            {7'd20,7'd46}:		p = 14'd920;
            {7'd20,7'd47}:		p = 14'd940;
            {7'd20,7'd48}:		p = 14'd960;
            {7'd20,7'd49}:		p = 14'd980;
            {7'd20,7'd50}:		p = 14'd1000;
            {7'd20,7'd51}:		p = 14'd1020;
            {7'd20,7'd52}:		p = 14'd1040;
            {7'd20,7'd53}:		p = 14'd1060;
            {7'd20,7'd54}:		p = 14'd1080;
            {7'd20,7'd55}:		p = 14'd1100;
            {7'd20,7'd56}:		p = 14'd1120;
            {7'd20,7'd57}:		p = 14'd1140;
            {7'd20,7'd58}:		p = 14'd1160;
            {7'd20,7'd59}:		p = 14'd1180;
            {7'd20,7'd60}:		p = 14'd1200;
            {7'd20,7'd61}:		p = 14'd1220;
            {7'd20,7'd62}:		p = 14'd1240;
            {7'd20,7'd63}:		p = 14'd1260;
            {7'd20,7'd64}:		p = 14'd1280;
            {7'd20,7'd65}:		p = 14'd1300;
            {7'd20,7'd66}:		p = 14'd1320;
            {7'd20,7'd67}:		p = 14'd1340;
            {7'd20,7'd68}:		p = 14'd1360;
            {7'd20,7'd69}:		p = 14'd1380;
            {7'd20,7'd70}:		p = 14'd1400;
            {7'd20,7'd71}:		p = 14'd1420;
            {7'd20,7'd72}:		p = 14'd1440;
            {7'd20,7'd73}:		p = 14'd1460;
            {7'd20,7'd74}:		p = 14'd1480;
            {7'd20,7'd75}:		p = 14'd1500;
            {7'd20,7'd76}:		p = 14'd1520;
            {7'd20,7'd77}:		p = 14'd1540;
            {7'd20,7'd78}:		p = 14'd1560;
            {7'd20,7'd79}:		p = 14'd1580;
            {7'd20,7'd80}:		p = 14'd1600;
            {7'd20,7'd81}:		p = 14'd1620;
            {7'd20,7'd82}:		p = 14'd1640;
            {7'd20,7'd83}:		p = 14'd1660;
            {7'd20,7'd84}:		p = 14'd1680;
            {7'd20,7'd85}:		p = 14'd1700;
            {7'd20,7'd86}:		p = 14'd1720;
            {7'd20,7'd87}:		p = 14'd1740;
            {7'd20,7'd88}:		p = 14'd1760;
            {7'd20,7'd89}:		p = 14'd1780;
            {7'd20,7'd90}:		p = 14'd1800;
            {7'd20,7'd91}:		p = 14'd1820;
            {7'd20,7'd92}:		p = 14'd1840;
            {7'd20,7'd93}:		p = 14'd1860;
            {7'd20,7'd94}:		p = 14'd1880;
            {7'd20,7'd95}:		p = 14'd1900;
            {7'd20,7'd96}:		p = 14'd1920;
            {7'd20,7'd97}:		p = 14'd1940;
            {7'd20,7'd98}:		p = 14'd1960;
            {7'd20,7'd99}:		p = 14'd1980;
            {7'd20,7'd100}:		p = 14'd2000;
            {7'd20,7'd101}:		p = 14'd2020;
            {7'd20,7'd102}:		p = 14'd2040;
            {7'd20,7'd103}:		p = 14'd2060;
            {7'd20,7'd104}:		p = 14'd2080;
            {7'd20,7'd105}:		p = 14'd2100;
            {7'd20,7'd106}:		p = 14'd2120;
            {7'd20,7'd107}:		p = 14'd2140;
            {7'd20,7'd108}:		p = 14'd2160;
            {7'd20,7'd109}:		p = 14'd2180;
            {7'd20,7'd110}:		p = 14'd2200;
            {7'd20,7'd111}:		p = 14'd2220;
            {7'd20,7'd112}:		p = 14'd2240;
            {7'd20,7'd113}:		p = 14'd2260;
            {7'd20,7'd114}:		p = 14'd2280;
            {7'd20,7'd115}:		p = 14'd2300;
            {7'd20,7'd116}:		p = 14'd2320;
            {7'd20,7'd117}:		p = 14'd2340;
            {7'd20,7'd118}:		p = 14'd2360;
            {7'd20,7'd119}:		p = 14'd2380;
            {7'd20,7'd120}:		p = 14'd2400;
            {7'd20,7'd121}:		p = 14'd2420;
            {7'd20,7'd122}:		p = 14'd2440;
            {7'd20,7'd123}:		p = 14'd2460;
            {7'd20,7'd124}:		p = 14'd2480;
            {7'd20,7'd125}:		p = 14'd2500;
            {7'd20,7'd126}:		p = 14'd2520;
            {7'd20,7'd127}:		p = 14'd2540;
            {7'd21,7'd0}:		p = 14'd0;
            {7'd21,7'd1}:		p = 14'd21;
            {7'd21,7'd2}:		p = 14'd42;
            {7'd21,7'd3}:		p = 14'd63;
            {7'd21,7'd4}:		p = 14'd84;
            {7'd21,7'd5}:		p = 14'd105;
            {7'd21,7'd6}:		p = 14'd126;
            {7'd21,7'd7}:		p = 14'd147;
            {7'd21,7'd8}:		p = 14'd168;
            {7'd21,7'd9}:		p = 14'd189;
            {7'd21,7'd10}:		p = 14'd210;
            {7'd21,7'd11}:		p = 14'd231;
            {7'd21,7'd12}:		p = 14'd252;
            {7'd21,7'd13}:		p = 14'd273;
            {7'd21,7'd14}:		p = 14'd294;
            {7'd21,7'd15}:		p = 14'd315;
            {7'd21,7'd16}:		p = 14'd336;
            {7'd21,7'd17}:		p = 14'd357;
            {7'd21,7'd18}:		p = 14'd378;
            {7'd21,7'd19}:		p = 14'd399;
            {7'd21,7'd20}:		p = 14'd420;
            {7'd21,7'd21}:		p = 14'd441;
            {7'd21,7'd22}:		p = 14'd462;
            {7'd21,7'd23}:		p = 14'd483;
            {7'd21,7'd24}:		p = 14'd504;
            {7'd21,7'd25}:		p = 14'd525;
            {7'd21,7'd26}:		p = 14'd546;
            {7'd21,7'd27}:		p = 14'd567;
            {7'd21,7'd28}:		p = 14'd588;
            {7'd21,7'd29}:		p = 14'd609;
            {7'd21,7'd30}:		p = 14'd630;
            {7'd21,7'd31}:		p = 14'd651;
            {7'd21,7'd32}:		p = 14'd672;
            {7'd21,7'd33}:		p = 14'd693;
            {7'd21,7'd34}:		p = 14'd714;
            {7'd21,7'd35}:		p = 14'd735;
            {7'd21,7'd36}:		p = 14'd756;
            {7'd21,7'd37}:		p = 14'd777;
            {7'd21,7'd38}:		p = 14'd798;
            {7'd21,7'd39}:		p = 14'd819;
            {7'd21,7'd40}:		p = 14'd840;
            {7'd21,7'd41}:		p = 14'd861;
            {7'd21,7'd42}:		p = 14'd882;
            {7'd21,7'd43}:		p = 14'd903;
            {7'd21,7'd44}:		p = 14'd924;
            {7'd21,7'd45}:		p = 14'd945;
            {7'd21,7'd46}:		p = 14'd966;
            {7'd21,7'd47}:		p = 14'd987;
            {7'd21,7'd48}:		p = 14'd1008;
            {7'd21,7'd49}:		p = 14'd1029;
            {7'd21,7'd50}:		p = 14'd1050;
            {7'd21,7'd51}:		p = 14'd1071;
            {7'd21,7'd52}:		p = 14'd1092;
            {7'd21,7'd53}:		p = 14'd1113;
            {7'd21,7'd54}:		p = 14'd1134;
            {7'd21,7'd55}:		p = 14'd1155;
            {7'd21,7'd56}:		p = 14'd1176;
            {7'd21,7'd57}:		p = 14'd1197;
            {7'd21,7'd58}:		p = 14'd1218;
            {7'd21,7'd59}:		p = 14'd1239;
            {7'd21,7'd60}:		p = 14'd1260;
            {7'd21,7'd61}:		p = 14'd1281;
            {7'd21,7'd62}:		p = 14'd1302;
            {7'd21,7'd63}:		p = 14'd1323;
            {7'd21,7'd64}:		p = 14'd1344;
            {7'd21,7'd65}:		p = 14'd1365;
            {7'd21,7'd66}:		p = 14'd1386;
            {7'd21,7'd67}:		p = 14'd1407;
            {7'd21,7'd68}:		p = 14'd1428;
            {7'd21,7'd69}:		p = 14'd1449;
            {7'd21,7'd70}:		p = 14'd1470;
            {7'd21,7'd71}:		p = 14'd1491;
            {7'd21,7'd72}:		p = 14'd1512;
            {7'd21,7'd73}:		p = 14'd1533;
            {7'd21,7'd74}:		p = 14'd1554;
            {7'd21,7'd75}:		p = 14'd1575;
            {7'd21,7'd76}:		p = 14'd1596;
            {7'd21,7'd77}:		p = 14'd1617;
            {7'd21,7'd78}:		p = 14'd1638;
            {7'd21,7'd79}:		p = 14'd1659;
            {7'd21,7'd80}:		p = 14'd1680;
            {7'd21,7'd81}:		p = 14'd1701;
            {7'd21,7'd82}:		p = 14'd1722;
            {7'd21,7'd83}:		p = 14'd1743;
            {7'd21,7'd84}:		p = 14'd1764;
            {7'd21,7'd85}:		p = 14'd1785;
            {7'd21,7'd86}:		p = 14'd1806;
            {7'd21,7'd87}:		p = 14'd1827;
            {7'd21,7'd88}:		p = 14'd1848;
            {7'd21,7'd89}:		p = 14'd1869;
            {7'd21,7'd90}:		p = 14'd1890;
            {7'd21,7'd91}:		p = 14'd1911;
            {7'd21,7'd92}:		p = 14'd1932;
            {7'd21,7'd93}:		p = 14'd1953;
            {7'd21,7'd94}:		p = 14'd1974;
            {7'd21,7'd95}:		p = 14'd1995;
            {7'd21,7'd96}:		p = 14'd2016;
            {7'd21,7'd97}:		p = 14'd2037;
            {7'd21,7'd98}:		p = 14'd2058;
            {7'd21,7'd99}:		p = 14'd2079;
            {7'd21,7'd100}:		p = 14'd2100;
            {7'd21,7'd101}:		p = 14'd2121;
            {7'd21,7'd102}:		p = 14'd2142;
            {7'd21,7'd103}:		p = 14'd2163;
            {7'd21,7'd104}:		p = 14'd2184;
            {7'd21,7'd105}:		p = 14'd2205;
            {7'd21,7'd106}:		p = 14'd2226;
            {7'd21,7'd107}:		p = 14'd2247;
            {7'd21,7'd108}:		p = 14'd2268;
            {7'd21,7'd109}:		p = 14'd2289;
            {7'd21,7'd110}:		p = 14'd2310;
            {7'd21,7'd111}:		p = 14'd2331;
            {7'd21,7'd112}:		p = 14'd2352;
            {7'd21,7'd113}:		p = 14'd2373;
            {7'd21,7'd114}:		p = 14'd2394;
            {7'd21,7'd115}:		p = 14'd2415;
            {7'd21,7'd116}:		p = 14'd2436;
            {7'd21,7'd117}:		p = 14'd2457;
            {7'd21,7'd118}:		p = 14'd2478;
            {7'd21,7'd119}:		p = 14'd2499;
            {7'd21,7'd120}:		p = 14'd2520;
            {7'd21,7'd121}:		p = 14'd2541;
            {7'd21,7'd122}:		p = 14'd2562;
            {7'd21,7'd123}:		p = 14'd2583;
            {7'd21,7'd124}:		p = 14'd2604;
            {7'd21,7'd125}:		p = 14'd2625;
            {7'd21,7'd126}:		p = 14'd2646;
            {7'd21,7'd127}:		p = 14'd2667;
            {7'd22,7'd0}:		p = 14'd0;
            {7'd22,7'd1}:		p = 14'd22;
            {7'd22,7'd2}:		p = 14'd44;
            {7'd22,7'd3}:		p = 14'd66;
            {7'd22,7'd4}:		p = 14'd88;
            {7'd22,7'd5}:		p = 14'd110;
            {7'd22,7'd6}:		p = 14'd132;
            {7'd22,7'd7}:		p = 14'd154;
            {7'd22,7'd8}:		p = 14'd176;
            {7'd22,7'd9}:		p = 14'd198;
            {7'd22,7'd10}:		p = 14'd220;
            {7'd22,7'd11}:		p = 14'd242;
            {7'd22,7'd12}:		p = 14'd264;
            {7'd22,7'd13}:		p = 14'd286;
            {7'd22,7'd14}:		p = 14'd308;
            {7'd22,7'd15}:		p = 14'd330;
            {7'd22,7'd16}:		p = 14'd352;
            {7'd22,7'd17}:		p = 14'd374;
            {7'd22,7'd18}:		p = 14'd396;
            {7'd22,7'd19}:		p = 14'd418;
            {7'd22,7'd20}:		p = 14'd440;
            {7'd22,7'd21}:		p = 14'd462;
            {7'd22,7'd22}:		p = 14'd484;
            {7'd22,7'd23}:		p = 14'd506;
            {7'd22,7'd24}:		p = 14'd528;
            {7'd22,7'd25}:		p = 14'd550;
            {7'd22,7'd26}:		p = 14'd572;
            {7'd22,7'd27}:		p = 14'd594;
            {7'd22,7'd28}:		p = 14'd616;
            {7'd22,7'd29}:		p = 14'd638;
            {7'd22,7'd30}:		p = 14'd660;
            {7'd22,7'd31}:		p = 14'd682;
            {7'd22,7'd32}:		p = 14'd704;
            {7'd22,7'd33}:		p = 14'd726;
            {7'd22,7'd34}:		p = 14'd748;
            {7'd22,7'd35}:		p = 14'd770;
            {7'd22,7'd36}:		p = 14'd792;
            {7'd22,7'd37}:		p = 14'd814;
            {7'd22,7'd38}:		p = 14'd836;
            {7'd22,7'd39}:		p = 14'd858;
            {7'd22,7'd40}:		p = 14'd880;
            {7'd22,7'd41}:		p = 14'd902;
            {7'd22,7'd42}:		p = 14'd924;
            {7'd22,7'd43}:		p = 14'd946;
            {7'd22,7'd44}:		p = 14'd968;
            {7'd22,7'd45}:		p = 14'd990;
            {7'd22,7'd46}:		p = 14'd1012;
            {7'd22,7'd47}:		p = 14'd1034;
            {7'd22,7'd48}:		p = 14'd1056;
            {7'd22,7'd49}:		p = 14'd1078;
            {7'd22,7'd50}:		p = 14'd1100;
            {7'd22,7'd51}:		p = 14'd1122;
            {7'd22,7'd52}:		p = 14'd1144;
            {7'd22,7'd53}:		p = 14'd1166;
            {7'd22,7'd54}:		p = 14'd1188;
            {7'd22,7'd55}:		p = 14'd1210;
            {7'd22,7'd56}:		p = 14'd1232;
            {7'd22,7'd57}:		p = 14'd1254;
            {7'd22,7'd58}:		p = 14'd1276;
            {7'd22,7'd59}:		p = 14'd1298;
            {7'd22,7'd60}:		p = 14'd1320;
            {7'd22,7'd61}:		p = 14'd1342;
            {7'd22,7'd62}:		p = 14'd1364;
            {7'd22,7'd63}:		p = 14'd1386;
            {7'd22,7'd64}:		p = 14'd1408;
            {7'd22,7'd65}:		p = 14'd1430;
            {7'd22,7'd66}:		p = 14'd1452;
            {7'd22,7'd67}:		p = 14'd1474;
            {7'd22,7'd68}:		p = 14'd1496;
            {7'd22,7'd69}:		p = 14'd1518;
            {7'd22,7'd70}:		p = 14'd1540;
            {7'd22,7'd71}:		p = 14'd1562;
            {7'd22,7'd72}:		p = 14'd1584;
            {7'd22,7'd73}:		p = 14'd1606;
            {7'd22,7'd74}:		p = 14'd1628;
            {7'd22,7'd75}:		p = 14'd1650;
            {7'd22,7'd76}:		p = 14'd1672;
            {7'd22,7'd77}:		p = 14'd1694;
            {7'd22,7'd78}:		p = 14'd1716;
            {7'd22,7'd79}:		p = 14'd1738;
            {7'd22,7'd80}:		p = 14'd1760;
            {7'd22,7'd81}:		p = 14'd1782;
            {7'd22,7'd82}:		p = 14'd1804;
            {7'd22,7'd83}:		p = 14'd1826;
            {7'd22,7'd84}:		p = 14'd1848;
            {7'd22,7'd85}:		p = 14'd1870;
            {7'd22,7'd86}:		p = 14'd1892;
            {7'd22,7'd87}:		p = 14'd1914;
            {7'd22,7'd88}:		p = 14'd1936;
            {7'd22,7'd89}:		p = 14'd1958;
            {7'd22,7'd90}:		p = 14'd1980;
            {7'd22,7'd91}:		p = 14'd2002;
            {7'd22,7'd92}:		p = 14'd2024;
            {7'd22,7'd93}:		p = 14'd2046;
            {7'd22,7'd94}:		p = 14'd2068;
            {7'd22,7'd95}:		p = 14'd2090;
            {7'd22,7'd96}:		p = 14'd2112;
            {7'd22,7'd97}:		p = 14'd2134;
            {7'd22,7'd98}:		p = 14'd2156;
            {7'd22,7'd99}:		p = 14'd2178;
            {7'd22,7'd100}:		p = 14'd2200;
            {7'd22,7'd101}:		p = 14'd2222;
            {7'd22,7'd102}:		p = 14'd2244;
            {7'd22,7'd103}:		p = 14'd2266;
            {7'd22,7'd104}:		p = 14'd2288;
            {7'd22,7'd105}:		p = 14'd2310;
            {7'd22,7'd106}:		p = 14'd2332;
            {7'd22,7'd107}:		p = 14'd2354;
            {7'd22,7'd108}:		p = 14'd2376;
            {7'd22,7'd109}:		p = 14'd2398;
            {7'd22,7'd110}:		p = 14'd2420;
            {7'd22,7'd111}:		p = 14'd2442;
            {7'd22,7'd112}:		p = 14'd2464;
            {7'd22,7'd113}:		p = 14'd2486;
            {7'd22,7'd114}:		p = 14'd2508;
            {7'd22,7'd115}:		p = 14'd2530;
            {7'd22,7'd116}:		p = 14'd2552;
            {7'd22,7'd117}:		p = 14'd2574;
            {7'd22,7'd118}:		p = 14'd2596;
            {7'd22,7'd119}:		p = 14'd2618;
            {7'd22,7'd120}:		p = 14'd2640;
            {7'd22,7'd121}:		p = 14'd2662;
            {7'd22,7'd122}:		p = 14'd2684;
            {7'd22,7'd123}:		p = 14'd2706;
            {7'd22,7'd124}:		p = 14'd2728;
            {7'd22,7'd125}:		p = 14'd2750;
            {7'd22,7'd126}:		p = 14'd2772;
            {7'd22,7'd127}:		p = 14'd2794;
            {7'd23,7'd0}:		p = 14'd0;
            {7'd23,7'd1}:		p = 14'd23;
            {7'd23,7'd2}:		p = 14'd46;
            {7'd23,7'd3}:		p = 14'd69;
            {7'd23,7'd4}:		p = 14'd92;
            {7'd23,7'd5}:		p = 14'd115;
            {7'd23,7'd6}:		p = 14'd138;
            {7'd23,7'd7}:		p = 14'd161;
            {7'd23,7'd8}:		p = 14'd184;
            {7'd23,7'd9}:		p = 14'd207;
            {7'd23,7'd10}:		p = 14'd230;
            {7'd23,7'd11}:		p = 14'd253;
            {7'd23,7'd12}:		p = 14'd276;
            {7'd23,7'd13}:		p = 14'd299;
            {7'd23,7'd14}:		p = 14'd322;
            {7'd23,7'd15}:		p = 14'd345;
            {7'd23,7'd16}:		p = 14'd368;
            {7'd23,7'd17}:		p = 14'd391;
            {7'd23,7'd18}:		p = 14'd414;
            {7'd23,7'd19}:		p = 14'd437;
            {7'd23,7'd20}:		p = 14'd460;
            {7'd23,7'd21}:		p = 14'd483;
            {7'd23,7'd22}:		p = 14'd506;
            {7'd23,7'd23}:		p = 14'd529;
            {7'd23,7'd24}:		p = 14'd552;
            {7'd23,7'd25}:		p = 14'd575;
            {7'd23,7'd26}:		p = 14'd598;
            {7'd23,7'd27}:		p = 14'd621;
            {7'd23,7'd28}:		p = 14'd644;
            {7'd23,7'd29}:		p = 14'd667;
            {7'd23,7'd30}:		p = 14'd690;
            {7'd23,7'd31}:		p = 14'd713;
            {7'd23,7'd32}:		p = 14'd736;
            {7'd23,7'd33}:		p = 14'd759;
            {7'd23,7'd34}:		p = 14'd782;
            {7'd23,7'd35}:		p = 14'd805;
            {7'd23,7'd36}:		p = 14'd828;
            {7'd23,7'd37}:		p = 14'd851;
            {7'd23,7'd38}:		p = 14'd874;
            {7'd23,7'd39}:		p = 14'd897;
            {7'd23,7'd40}:		p = 14'd920;
            {7'd23,7'd41}:		p = 14'd943;
            {7'd23,7'd42}:		p = 14'd966;
            {7'd23,7'd43}:		p = 14'd989;
            {7'd23,7'd44}:		p = 14'd1012;
            {7'd23,7'd45}:		p = 14'd1035;
            {7'd23,7'd46}:		p = 14'd1058;
            {7'd23,7'd47}:		p = 14'd1081;
            {7'd23,7'd48}:		p = 14'd1104;
            {7'd23,7'd49}:		p = 14'd1127;
            {7'd23,7'd50}:		p = 14'd1150;
            {7'd23,7'd51}:		p = 14'd1173;
            {7'd23,7'd52}:		p = 14'd1196;
            {7'd23,7'd53}:		p = 14'd1219;
            {7'd23,7'd54}:		p = 14'd1242;
            {7'd23,7'd55}:		p = 14'd1265;
            {7'd23,7'd56}:		p = 14'd1288;
            {7'd23,7'd57}:		p = 14'd1311;
            {7'd23,7'd58}:		p = 14'd1334;
            {7'd23,7'd59}:		p = 14'd1357;
            {7'd23,7'd60}:		p = 14'd1380;
            {7'd23,7'd61}:		p = 14'd1403;
            {7'd23,7'd62}:		p = 14'd1426;
            {7'd23,7'd63}:		p = 14'd1449;
            {7'd23,7'd64}:		p = 14'd1472;
            {7'd23,7'd65}:		p = 14'd1495;
            {7'd23,7'd66}:		p = 14'd1518;
            {7'd23,7'd67}:		p = 14'd1541;
            {7'd23,7'd68}:		p = 14'd1564;
            {7'd23,7'd69}:		p = 14'd1587;
            {7'd23,7'd70}:		p = 14'd1610;
            {7'd23,7'd71}:		p = 14'd1633;
            {7'd23,7'd72}:		p = 14'd1656;
            {7'd23,7'd73}:		p = 14'd1679;
            {7'd23,7'd74}:		p = 14'd1702;
            {7'd23,7'd75}:		p = 14'd1725;
            {7'd23,7'd76}:		p = 14'd1748;
            {7'd23,7'd77}:		p = 14'd1771;
            {7'd23,7'd78}:		p = 14'd1794;
            {7'd23,7'd79}:		p = 14'd1817;
            {7'd23,7'd80}:		p = 14'd1840;
            {7'd23,7'd81}:		p = 14'd1863;
            {7'd23,7'd82}:		p = 14'd1886;
            {7'd23,7'd83}:		p = 14'd1909;
            {7'd23,7'd84}:		p = 14'd1932;
            {7'd23,7'd85}:		p = 14'd1955;
            {7'd23,7'd86}:		p = 14'd1978;
            {7'd23,7'd87}:		p = 14'd2001;
            {7'd23,7'd88}:		p = 14'd2024;
            {7'd23,7'd89}:		p = 14'd2047;
            {7'd23,7'd90}:		p = 14'd2070;
            {7'd23,7'd91}:		p = 14'd2093;
            {7'd23,7'd92}:		p = 14'd2116;
            {7'd23,7'd93}:		p = 14'd2139;
            {7'd23,7'd94}:		p = 14'd2162;
            {7'd23,7'd95}:		p = 14'd2185;
            {7'd23,7'd96}:		p = 14'd2208;
            {7'd23,7'd97}:		p = 14'd2231;
            {7'd23,7'd98}:		p = 14'd2254;
            {7'd23,7'd99}:		p = 14'd2277;
            {7'd23,7'd100}:		p = 14'd2300;
            {7'd23,7'd101}:		p = 14'd2323;
            {7'd23,7'd102}:		p = 14'd2346;
            {7'd23,7'd103}:		p = 14'd2369;
            {7'd23,7'd104}:		p = 14'd2392;
            {7'd23,7'd105}:		p = 14'd2415;
            {7'd23,7'd106}:		p = 14'd2438;
            {7'd23,7'd107}:		p = 14'd2461;
            {7'd23,7'd108}:		p = 14'd2484;
            {7'd23,7'd109}:		p = 14'd2507;
            {7'd23,7'd110}:		p = 14'd2530;
            {7'd23,7'd111}:		p = 14'd2553;
            {7'd23,7'd112}:		p = 14'd2576;
            {7'd23,7'd113}:		p = 14'd2599;
            {7'd23,7'd114}:		p = 14'd2622;
            {7'd23,7'd115}:		p = 14'd2645;
            {7'd23,7'd116}:		p = 14'd2668;
            {7'd23,7'd117}:		p = 14'd2691;
            {7'd23,7'd118}:		p = 14'd2714;
            {7'd23,7'd119}:		p = 14'd2737;
            {7'd23,7'd120}:		p = 14'd2760;
            {7'd23,7'd121}:		p = 14'd2783;
            {7'd23,7'd122}:		p = 14'd2806;
            {7'd23,7'd123}:		p = 14'd2829;
            {7'd23,7'd124}:		p = 14'd2852;
            {7'd23,7'd125}:		p = 14'd2875;
            {7'd23,7'd126}:		p = 14'd2898;
            {7'd23,7'd127}:		p = 14'd2921;
            {7'd24,7'd0}:		p = 14'd0;
            {7'd24,7'd1}:		p = 14'd24;
            {7'd24,7'd2}:		p = 14'd48;
            {7'd24,7'd3}:		p = 14'd72;
            {7'd24,7'd4}:		p = 14'd96;
            {7'd24,7'd5}:		p = 14'd120;
            {7'd24,7'd6}:		p = 14'd144;
            {7'd24,7'd7}:		p = 14'd168;
            {7'd24,7'd8}:		p = 14'd192;
            {7'd24,7'd9}:		p = 14'd216;
            {7'd24,7'd10}:		p = 14'd240;
            {7'd24,7'd11}:		p = 14'd264;
            {7'd24,7'd12}:		p = 14'd288;
            {7'd24,7'd13}:		p = 14'd312;
            {7'd24,7'd14}:		p = 14'd336;
            {7'd24,7'd15}:		p = 14'd360;
            {7'd24,7'd16}:		p = 14'd384;
            {7'd24,7'd17}:		p = 14'd408;
            {7'd24,7'd18}:		p = 14'd432;
            {7'd24,7'd19}:		p = 14'd456;
            {7'd24,7'd20}:		p = 14'd480;
            {7'd24,7'd21}:		p = 14'd504;
            {7'd24,7'd22}:		p = 14'd528;
            {7'd24,7'd23}:		p = 14'd552;
            {7'd24,7'd24}:		p = 14'd576;
            {7'd24,7'd25}:		p = 14'd600;
            {7'd24,7'd26}:		p = 14'd624;
            {7'd24,7'd27}:		p = 14'd648;
            {7'd24,7'd28}:		p = 14'd672;
            {7'd24,7'd29}:		p = 14'd696;
            {7'd24,7'd30}:		p = 14'd720;
            {7'd24,7'd31}:		p = 14'd744;
            {7'd24,7'd32}:		p = 14'd768;
            {7'd24,7'd33}:		p = 14'd792;
            {7'd24,7'd34}:		p = 14'd816;
            {7'd24,7'd35}:		p = 14'd840;
            {7'd24,7'd36}:		p = 14'd864;
            {7'd24,7'd37}:		p = 14'd888;
            {7'd24,7'd38}:		p = 14'd912;
            {7'd24,7'd39}:		p = 14'd936;
            {7'd24,7'd40}:		p = 14'd960;
            {7'd24,7'd41}:		p = 14'd984;
            {7'd24,7'd42}:		p = 14'd1008;
            {7'd24,7'd43}:		p = 14'd1032;
            {7'd24,7'd44}:		p = 14'd1056;
            {7'd24,7'd45}:		p = 14'd1080;
            {7'd24,7'd46}:		p = 14'd1104;
            {7'd24,7'd47}:		p = 14'd1128;
            {7'd24,7'd48}:		p = 14'd1152;
            {7'd24,7'd49}:		p = 14'd1176;
            {7'd24,7'd50}:		p = 14'd1200;
            {7'd24,7'd51}:		p = 14'd1224;
            {7'd24,7'd52}:		p = 14'd1248;
            {7'd24,7'd53}:		p = 14'd1272;
            {7'd24,7'd54}:		p = 14'd1296;
            {7'd24,7'd55}:		p = 14'd1320;
            {7'd24,7'd56}:		p = 14'd1344;
            {7'd24,7'd57}:		p = 14'd1368;
            {7'd24,7'd58}:		p = 14'd1392;
            {7'd24,7'd59}:		p = 14'd1416;
            {7'd24,7'd60}:		p = 14'd1440;
            {7'd24,7'd61}:		p = 14'd1464;
            {7'd24,7'd62}:		p = 14'd1488;
            {7'd24,7'd63}:		p = 14'd1512;
            {7'd24,7'd64}:		p = 14'd1536;
            {7'd24,7'd65}:		p = 14'd1560;
            {7'd24,7'd66}:		p = 14'd1584;
            {7'd24,7'd67}:		p = 14'd1608;
            {7'd24,7'd68}:		p = 14'd1632;
            {7'd24,7'd69}:		p = 14'd1656;
            {7'd24,7'd70}:		p = 14'd1680;
            {7'd24,7'd71}:		p = 14'd1704;
            {7'd24,7'd72}:		p = 14'd1728;
            {7'd24,7'd73}:		p = 14'd1752;
            {7'd24,7'd74}:		p = 14'd1776;
            {7'd24,7'd75}:		p = 14'd1800;
            {7'd24,7'd76}:		p = 14'd1824;
            {7'd24,7'd77}:		p = 14'd1848;
            {7'd24,7'd78}:		p = 14'd1872;
            {7'd24,7'd79}:		p = 14'd1896;
            {7'd24,7'd80}:		p = 14'd1920;
            {7'd24,7'd81}:		p = 14'd1944;
            {7'd24,7'd82}:		p = 14'd1968;
            {7'd24,7'd83}:		p = 14'd1992;
            {7'd24,7'd84}:		p = 14'd2016;
            {7'd24,7'd85}:		p = 14'd2040;
            {7'd24,7'd86}:		p = 14'd2064;
            {7'd24,7'd87}:		p = 14'd2088;
            {7'd24,7'd88}:		p = 14'd2112;
            {7'd24,7'd89}:		p = 14'd2136;
            {7'd24,7'd90}:		p = 14'd2160;
            {7'd24,7'd91}:		p = 14'd2184;
            {7'd24,7'd92}:		p = 14'd2208;
            {7'd24,7'd93}:		p = 14'd2232;
            {7'd24,7'd94}:		p = 14'd2256;
            {7'd24,7'd95}:		p = 14'd2280;
            {7'd24,7'd96}:		p = 14'd2304;
            {7'd24,7'd97}:		p = 14'd2328;
            {7'd24,7'd98}:		p = 14'd2352;
            {7'd24,7'd99}:		p = 14'd2376;
            {7'd24,7'd100}:		p = 14'd2400;
            {7'd24,7'd101}:		p = 14'd2424;
            {7'd24,7'd102}:		p = 14'd2448;
            {7'd24,7'd103}:		p = 14'd2472;
            {7'd24,7'd104}:		p = 14'd2496;
            {7'd24,7'd105}:		p = 14'd2520;
            {7'd24,7'd106}:		p = 14'd2544;
            {7'd24,7'd107}:		p = 14'd2568;
            {7'd24,7'd108}:		p = 14'd2592;
            {7'd24,7'd109}:		p = 14'd2616;
            {7'd24,7'd110}:		p = 14'd2640;
            {7'd24,7'd111}:		p = 14'd2664;
            {7'd24,7'd112}:		p = 14'd2688;
            {7'd24,7'd113}:		p = 14'd2712;
            {7'd24,7'd114}:		p = 14'd2736;
            {7'd24,7'd115}:		p = 14'd2760;
            {7'd24,7'd116}:		p = 14'd2784;
            {7'd24,7'd117}:		p = 14'd2808;
            {7'd24,7'd118}:		p = 14'd2832;
            {7'd24,7'd119}:		p = 14'd2856;
            {7'd24,7'd120}:		p = 14'd2880;
            {7'd24,7'd121}:		p = 14'd2904;
            {7'd24,7'd122}:		p = 14'd2928;
            {7'd24,7'd123}:		p = 14'd2952;
            {7'd24,7'd124}:		p = 14'd2976;
            {7'd24,7'd125}:		p = 14'd3000;
            {7'd24,7'd126}:		p = 14'd3024;
            {7'd24,7'd127}:		p = 14'd3048;
            {7'd25,7'd0}:		p = 14'd0;
            {7'd25,7'd1}:		p = 14'd25;
            {7'd25,7'd2}:		p = 14'd50;
            {7'd25,7'd3}:		p = 14'd75;
            {7'd25,7'd4}:		p = 14'd100;
            {7'd25,7'd5}:		p = 14'd125;
            {7'd25,7'd6}:		p = 14'd150;
            {7'd25,7'd7}:		p = 14'd175;
            {7'd25,7'd8}:		p = 14'd200;
            {7'd25,7'd9}:		p = 14'd225;
            {7'd25,7'd10}:		p = 14'd250;
            {7'd25,7'd11}:		p = 14'd275;
            {7'd25,7'd12}:		p = 14'd300;
            {7'd25,7'd13}:		p = 14'd325;
            {7'd25,7'd14}:		p = 14'd350;
            {7'd25,7'd15}:		p = 14'd375;
            {7'd25,7'd16}:		p = 14'd400;
            {7'd25,7'd17}:		p = 14'd425;
            {7'd25,7'd18}:		p = 14'd450;
            {7'd25,7'd19}:		p = 14'd475;
            {7'd25,7'd20}:		p = 14'd500;
            {7'd25,7'd21}:		p = 14'd525;
            {7'd25,7'd22}:		p = 14'd550;
            {7'd25,7'd23}:		p = 14'd575;
            {7'd25,7'd24}:		p = 14'd600;
            {7'd25,7'd25}:		p = 14'd625;
            {7'd25,7'd26}:		p = 14'd650;
            {7'd25,7'd27}:		p = 14'd675;
            {7'd25,7'd28}:		p = 14'd700;
            {7'd25,7'd29}:		p = 14'd725;
            {7'd25,7'd30}:		p = 14'd750;
            {7'd25,7'd31}:		p = 14'd775;
            {7'd25,7'd32}:		p = 14'd800;
            {7'd25,7'd33}:		p = 14'd825;
            {7'd25,7'd34}:		p = 14'd850;
            {7'd25,7'd35}:		p = 14'd875;
            {7'd25,7'd36}:		p = 14'd900;
            {7'd25,7'd37}:		p = 14'd925;
            {7'd25,7'd38}:		p = 14'd950;
            {7'd25,7'd39}:		p = 14'd975;
            {7'd25,7'd40}:		p = 14'd1000;
            {7'd25,7'd41}:		p = 14'd1025;
            {7'd25,7'd42}:		p = 14'd1050;
            {7'd25,7'd43}:		p = 14'd1075;
            {7'd25,7'd44}:		p = 14'd1100;
            {7'd25,7'd45}:		p = 14'd1125;
            {7'd25,7'd46}:		p = 14'd1150;
            {7'd25,7'd47}:		p = 14'd1175;
            {7'd25,7'd48}:		p = 14'd1200;
            {7'd25,7'd49}:		p = 14'd1225;
            {7'd25,7'd50}:		p = 14'd1250;
            {7'd25,7'd51}:		p = 14'd1275;
            {7'd25,7'd52}:		p = 14'd1300;
            {7'd25,7'd53}:		p = 14'd1325;
            {7'd25,7'd54}:		p = 14'd1350;
            {7'd25,7'd55}:		p = 14'd1375;
            {7'd25,7'd56}:		p = 14'd1400;
            {7'd25,7'd57}:		p = 14'd1425;
            {7'd25,7'd58}:		p = 14'd1450;
            {7'd25,7'd59}:		p = 14'd1475;
            {7'd25,7'd60}:		p = 14'd1500;
            {7'd25,7'd61}:		p = 14'd1525;
            {7'd25,7'd62}:		p = 14'd1550;
            {7'd25,7'd63}:		p = 14'd1575;
            {7'd25,7'd64}:		p = 14'd1600;
            {7'd25,7'd65}:		p = 14'd1625;
            {7'd25,7'd66}:		p = 14'd1650;
            {7'd25,7'd67}:		p = 14'd1675;
            {7'd25,7'd68}:		p = 14'd1700;
            {7'd25,7'd69}:		p = 14'd1725;
            {7'd25,7'd70}:		p = 14'd1750;
            {7'd25,7'd71}:		p = 14'd1775;
            {7'd25,7'd72}:		p = 14'd1800;
            {7'd25,7'd73}:		p = 14'd1825;
            {7'd25,7'd74}:		p = 14'd1850;
            {7'd25,7'd75}:		p = 14'd1875;
            {7'd25,7'd76}:		p = 14'd1900;
            {7'd25,7'd77}:		p = 14'd1925;
            {7'd25,7'd78}:		p = 14'd1950;
            {7'd25,7'd79}:		p = 14'd1975;
            {7'd25,7'd80}:		p = 14'd2000;
            {7'd25,7'd81}:		p = 14'd2025;
            {7'd25,7'd82}:		p = 14'd2050;
            {7'd25,7'd83}:		p = 14'd2075;
            {7'd25,7'd84}:		p = 14'd2100;
            {7'd25,7'd85}:		p = 14'd2125;
            {7'd25,7'd86}:		p = 14'd2150;
            {7'd25,7'd87}:		p = 14'd2175;
            {7'd25,7'd88}:		p = 14'd2200;
            {7'd25,7'd89}:		p = 14'd2225;
            {7'd25,7'd90}:		p = 14'd2250;
            {7'd25,7'd91}:		p = 14'd2275;
            {7'd25,7'd92}:		p = 14'd2300;
            {7'd25,7'd93}:		p = 14'd2325;
            {7'd25,7'd94}:		p = 14'd2350;
            {7'd25,7'd95}:		p = 14'd2375;
            {7'd25,7'd96}:		p = 14'd2400;
            {7'd25,7'd97}:		p = 14'd2425;
            {7'd25,7'd98}:		p = 14'd2450;
            {7'd25,7'd99}:		p = 14'd2475;
            {7'd25,7'd100}:		p = 14'd2500;
            {7'd25,7'd101}:		p = 14'd2525;
            {7'd25,7'd102}:		p = 14'd2550;
            {7'd25,7'd103}:		p = 14'd2575;
            {7'd25,7'd104}:		p = 14'd2600;
            {7'd25,7'd105}:		p = 14'd2625;
            {7'd25,7'd106}:		p = 14'd2650;
            {7'd25,7'd107}:		p = 14'd2675;
            {7'd25,7'd108}:		p = 14'd2700;
            {7'd25,7'd109}:		p = 14'd2725;
            {7'd25,7'd110}:		p = 14'd2750;
            {7'd25,7'd111}:		p = 14'd2775;
            {7'd25,7'd112}:		p = 14'd2800;
            {7'd25,7'd113}:		p = 14'd2825;
            {7'd25,7'd114}:		p = 14'd2850;
            {7'd25,7'd115}:		p = 14'd2875;
            {7'd25,7'd116}:		p = 14'd2900;
            {7'd25,7'd117}:		p = 14'd2925;
            {7'd25,7'd118}:		p = 14'd2950;
            {7'd25,7'd119}:		p = 14'd2975;
            {7'd25,7'd120}:		p = 14'd3000;
            {7'd25,7'd121}:		p = 14'd3025;
            {7'd25,7'd122}:		p = 14'd3050;
            {7'd25,7'd123}:		p = 14'd3075;
            {7'd25,7'd124}:		p = 14'd3100;
            {7'd25,7'd125}:		p = 14'd3125;
            {7'd25,7'd126}:		p = 14'd3150;
            {7'd25,7'd127}:		p = 14'd3175;
            {7'd26,7'd0}:		p = 14'd0;
            {7'd26,7'd1}:		p = 14'd26;
            {7'd26,7'd2}:		p = 14'd52;
            {7'd26,7'd3}:		p = 14'd78;
            {7'd26,7'd4}:		p = 14'd104;
            {7'd26,7'd5}:		p = 14'd130;
            {7'd26,7'd6}:		p = 14'd156;
            {7'd26,7'd7}:		p = 14'd182;
            {7'd26,7'd8}:		p = 14'd208;
            {7'd26,7'd9}:		p = 14'd234;
            {7'd26,7'd10}:		p = 14'd260;
            {7'd26,7'd11}:		p = 14'd286;
            {7'd26,7'd12}:		p = 14'd312;
            {7'd26,7'd13}:		p = 14'd338;
            {7'd26,7'd14}:		p = 14'd364;
            {7'd26,7'd15}:		p = 14'd390;
            {7'd26,7'd16}:		p = 14'd416;
            {7'd26,7'd17}:		p = 14'd442;
            {7'd26,7'd18}:		p = 14'd468;
            {7'd26,7'd19}:		p = 14'd494;
            {7'd26,7'd20}:		p = 14'd520;
            {7'd26,7'd21}:		p = 14'd546;
            {7'd26,7'd22}:		p = 14'd572;
            {7'd26,7'd23}:		p = 14'd598;
            {7'd26,7'd24}:		p = 14'd624;
            {7'd26,7'd25}:		p = 14'd650;
            {7'd26,7'd26}:		p = 14'd676;
            {7'd26,7'd27}:		p = 14'd702;
            {7'd26,7'd28}:		p = 14'd728;
            {7'd26,7'd29}:		p = 14'd754;
            {7'd26,7'd30}:		p = 14'd780;
            {7'd26,7'd31}:		p = 14'd806;
            {7'd26,7'd32}:		p = 14'd832;
            {7'd26,7'd33}:		p = 14'd858;
            {7'd26,7'd34}:		p = 14'd884;
            {7'd26,7'd35}:		p = 14'd910;
            {7'd26,7'd36}:		p = 14'd936;
            {7'd26,7'd37}:		p = 14'd962;
            {7'd26,7'd38}:		p = 14'd988;
            {7'd26,7'd39}:		p = 14'd1014;
            {7'd26,7'd40}:		p = 14'd1040;
            {7'd26,7'd41}:		p = 14'd1066;
            {7'd26,7'd42}:		p = 14'd1092;
            {7'd26,7'd43}:		p = 14'd1118;
            {7'd26,7'd44}:		p = 14'd1144;
            {7'd26,7'd45}:		p = 14'd1170;
            {7'd26,7'd46}:		p = 14'd1196;
            {7'd26,7'd47}:		p = 14'd1222;
            {7'd26,7'd48}:		p = 14'd1248;
            {7'd26,7'd49}:		p = 14'd1274;
            {7'd26,7'd50}:		p = 14'd1300;
            {7'd26,7'd51}:		p = 14'd1326;
            {7'd26,7'd52}:		p = 14'd1352;
            {7'd26,7'd53}:		p = 14'd1378;
            {7'd26,7'd54}:		p = 14'd1404;
            {7'd26,7'd55}:		p = 14'd1430;
            {7'd26,7'd56}:		p = 14'd1456;
            {7'd26,7'd57}:		p = 14'd1482;
            {7'd26,7'd58}:		p = 14'd1508;
            {7'd26,7'd59}:		p = 14'd1534;
            {7'd26,7'd60}:		p = 14'd1560;
            {7'd26,7'd61}:		p = 14'd1586;
            {7'd26,7'd62}:		p = 14'd1612;
            {7'd26,7'd63}:		p = 14'd1638;
            {7'd26,7'd64}:		p = 14'd1664;
            {7'd26,7'd65}:		p = 14'd1690;
            {7'd26,7'd66}:		p = 14'd1716;
            {7'd26,7'd67}:		p = 14'd1742;
            {7'd26,7'd68}:		p = 14'd1768;
            {7'd26,7'd69}:		p = 14'd1794;
            {7'd26,7'd70}:		p = 14'd1820;
            {7'd26,7'd71}:		p = 14'd1846;
            {7'd26,7'd72}:		p = 14'd1872;
            {7'd26,7'd73}:		p = 14'd1898;
            {7'd26,7'd74}:		p = 14'd1924;
            {7'd26,7'd75}:		p = 14'd1950;
            {7'd26,7'd76}:		p = 14'd1976;
            {7'd26,7'd77}:		p = 14'd2002;
            {7'd26,7'd78}:		p = 14'd2028;
            {7'd26,7'd79}:		p = 14'd2054;
            {7'd26,7'd80}:		p = 14'd2080;
            {7'd26,7'd81}:		p = 14'd2106;
            {7'd26,7'd82}:		p = 14'd2132;
            {7'd26,7'd83}:		p = 14'd2158;
            {7'd26,7'd84}:		p = 14'd2184;
            {7'd26,7'd85}:		p = 14'd2210;
            {7'd26,7'd86}:		p = 14'd2236;
            {7'd26,7'd87}:		p = 14'd2262;
            {7'd26,7'd88}:		p = 14'd2288;
            {7'd26,7'd89}:		p = 14'd2314;
            {7'd26,7'd90}:		p = 14'd2340;
            {7'd26,7'd91}:		p = 14'd2366;
            {7'd26,7'd92}:		p = 14'd2392;
            {7'd26,7'd93}:		p = 14'd2418;
            {7'd26,7'd94}:		p = 14'd2444;
            {7'd26,7'd95}:		p = 14'd2470;
            {7'd26,7'd96}:		p = 14'd2496;
            {7'd26,7'd97}:		p = 14'd2522;
            {7'd26,7'd98}:		p = 14'd2548;
            {7'd26,7'd99}:		p = 14'd2574;
            {7'd26,7'd100}:		p = 14'd2600;
            {7'd26,7'd101}:		p = 14'd2626;
            {7'd26,7'd102}:		p = 14'd2652;
            {7'd26,7'd103}:		p = 14'd2678;
            {7'd26,7'd104}:		p = 14'd2704;
            {7'd26,7'd105}:		p = 14'd2730;
            {7'd26,7'd106}:		p = 14'd2756;
            {7'd26,7'd107}:		p = 14'd2782;
            {7'd26,7'd108}:		p = 14'd2808;
            {7'd26,7'd109}:		p = 14'd2834;
            {7'd26,7'd110}:		p = 14'd2860;
            {7'd26,7'd111}:		p = 14'd2886;
            {7'd26,7'd112}:		p = 14'd2912;
            {7'd26,7'd113}:		p = 14'd2938;
            {7'd26,7'd114}:		p = 14'd2964;
            {7'd26,7'd115}:		p = 14'd2990;
            {7'd26,7'd116}:		p = 14'd3016;
            {7'd26,7'd117}:		p = 14'd3042;
            {7'd26,7'd118}:		p = 14'd3068;
            {7'd26,7'd119}:		p = 14'd3094;
            {7'd26,7'd120}:		p = 14'd3120;
            {7'd26,7'd121}:		p = 14'd3146;
            {7'd26,7'd122}:		p = 14'd3172;
            {7'd26,7'd123}:		p = 14'd3198;
            {7'd26,7'd124}:		p = 14'd3224;
            {7'd26,7'd125}:		p = 14'd3250;
            {7'd26,7'd126}:		p = 14'd3276;
            {7'd26,7'd127}:		p = 14'd3302;
            {7'd27,7'd0}:		p = 14'd0;
            {7'd27,7'd1}:		p = 14'd27;
            {7'd27,7'd2}:		p = 14'd54;
            {7'd27,7'd3}:		p = 14'd81;
            {7'd27,7'd4}:		p = 14'd108;
            {7'd27,7'd5}:		p = 14'd135;
            {7'd27,7'd6}:		p = 14'd162;
            {7'd27,7'd7}:		p = 14'd189;
            {7'd27,7'd8}:		p = 14'd216;
            {7'd27,7'd9}:		p = 14'd243;
            {7'd27,7'd10}:		p = 14'd270;
            {7'd27,7'd11}:		p = 14'd297;
            {7'd27,7'd12}:		p = 14'd324;
            {7'd27,7'd13}:		p = 14'd351;
            {7'd27,7'd14}:		p = 14'd378;
            {7'd27,7'd15}:		p = 14'd405;
            {7'd27,7'd16}:		p = 14'd432;
            {7'd27,7'd17}:		p = 14'd459;
            {7'd27,7'd18}:		p = 14'd486;
            {7'd27,7'd19}:		p = 14'd513;
            {7'd27,7'd20}:		p = 14'd540;
            {7'd27,7'd21}:		p = 14'd567;
            {7'd27,7'd22}:		p = 14'd594;
            {7'd27,7'd23}:		p = 14'd621;
            {7'd27,7'd24}:		p = 14'd648;
            {7'd27,7'd25}:		p = 14'd675;
            {7'd27,7'd26}:		p = 14'd702;
            {7'd27,7'd27}:		p = 14'd729;
            {7'd27,7'd28}:		p = 14'd756;
            {7'd27,7'd29}:		p = 14'd783;
            {7'd27,7'd30}:		p = 14'd810;
            {7'd27,7'd31}:		p = 14'd837;
            {7'd27,7'd32}:		p = 14'd864;
            {7'd27,7'd33}:		p = 14'd891;
            {7'd27,7'd34}:		p = 14'd918;
            {7'd27,7'd35}:		p = 14'd945;
            {7'd27,7'd36}:		p = 14'd972;
            {7'd27,7'd37}:		p = 14'd999;
            {7'd27,7'd38}:		p = 14'd1026;
            {7'd27,7'd39}:		p = 14'd1053;
            {7'd27,7'd40}:		p = 14'd1080;
            {7'd27,7'd41}:		p = 14'd1107;
            {7'd27,7'd42}:		p = 14'd1134;
            {7'd27,7'd43}:		p = 14'd1161;
            {7'd27,7'd44}:		p = 14'd1188;
            {7'd27,7'd45}:		p = 14'd1215;
            {7'd27,7'd46}:		p = 14'd1242;
            {7'd27,7'd47}:		p = 14'd1269;
            {7'd27,7'd48}:		p = 14'd1296;
            {7'd27,7'd49}:		p = 14'd1323;
            {7'd27,7'd50}:		p = 14'd1350;
            {7'd27,7'd51}:		p = 14'd1377;
            {7'd27,7'd52}:		p = 14'd1404;
            {7'd27,7'd53}:		p = 14'd1431;
            {7'd27,7'd54}:		p = 14'd1458;
            {7'd27,7'd55}:		p = 14'd1485;
            {7'd27,7'd56}:		p = 14'd1512;
            {7'd27,7'd57}:		p = 14'd1539;
            {7'd27,7'd58}:		p = 14'd1566;
            {7'd27,7'd59}:		p = 14'd1593;
            {7'd27,7'd60}:		p = 14'd1620;
            {7'd27,7'd61}:		p = 14'd1647;
            {7'd27,7'd62}:		p = 14'd1674;
            {7'd27,7'd63}:		p = 14'd1701;
            {7'd27,7'd64}:		p = 14'd1728;
            {7'd27,7'd65}:		p = 14'd1755;
            {7'd27,7'd66}:		p = 14'd1782;
            {7'd27,7'd67}:		p = 14'd1809;
            {7'd27,7'd68}:		p = 14'd1836;
            {7'd27,7'd69}:		p = 14'd1863;
            {7'd27,7'd70}:		p = 14'd1890;
            {7'd27,7'd71}:		p = 14'd1917;
            {7'd27,7'd72}:		p = 14'd1944;
            {7'd27,7'd73}:		p = 14'd1971;
            {7'd27,7'd74}:		p = 14'd1998;
            {7'd27,7'd75}:		p = 14'd2025;
            {7'd27,7'd76}:		p = 14'd2052;
            {7'd27,7'd77}:		p = 14'd2079;
            {7'd27,7'd78}:		p = 14'd2106;
            {7'd27,7'd79}:		p = 14'd2133;
            {7'd27,7'd80}:		p = 14'd2160;
            {7'd27,7'd81}:		p = 14'd2187;
            {7'd27,7'd82}:		p = 14'd2214;
            {7'd27,7'd83}:		p = 14'd2241;
            {7'd27,7'd84}:		p = 14'd2268;
            {7'd27,7'd85}:		p = 14'd2295;
            {7'd27,7'd86}:		p = 14'd2322;
            {7'd27,7'd87}:		p = 14'd2349;
            {7'd27,7'd88}:		p = 14'd2376;
            {7'd27,7'd89}:		p = 14'd2403;
            {7'd27,7'd90}:		p = 14'd2430;
            {7'd27,7'd91}:		p = 14'd2457;
            {7'd27,7'd92}:		p = 14'd2484;
            {7'd27,7'd93}:		p = 14'd2511;
            {7'd27,7'd94}:		p = 14'd2538;
            {7'd27,7'd95}:		p = 14'd2565;
            {7'd27,7'd96}:		p = 14'd2592;
            {7'd27,7'd97}:		p = 14'd2619;
            {7'd27,7'd98}:		p = 14'd2646;
            {7'd27,7'd99}:		p = 14'd2673;
            {7'd27,7'd100}:		p = 14'd2700;
            {7'd27,7'd101}:		p = 14'd2727;
            {7'd27,7'd102}:		p = 14'd2754;
            {7'd27,7'd103}:		p = 14'd2781;
            {7'd27,7'd104}:		p = 14'd2808;
            {7'd27,7'd105}:		p = 14'd2835;
            {7'd27,7'd106}:		p = 14'd2862;
            {7'd27,7'd107}:		p = 14'd2889;
            {7'd27,7'd108}:		p = 14'd2916;
            {7'd27,7'd109}:		p = 14'd2943;
            {7'd27,7'd110}:		p = 14'd2970;
            {7'd27,7'd111}:		p = 14'd2997;
            {7'd27,7'd112}:		p = 14'd3024;
            {7'd27,7'd113}:		p = 14'd3051;
            {7'd27,7'd114}:		p = 14'd3078;
            {7'd27,7'd115}:		p = 14'd3105;
            {7'd27,7'd116}:		p = 14'd3132;
            {7'd27,7'd117}:		p = 14'd3159;
            {7'd27,7'd118}:		p = 14'd3186;
            {7'd27,7'd119}:		p = 14'd3213;
            {7'd27,7'd120}:		p = 14'd3240;
            {7'd27,7'd121}:		p = 14'd3267;
            {7'd27,7'd122}:		p = 14'd3294;
            {7'd27,7'd123}:		p = 14'd3321;
            {7'd27,7'd124}:		p = 14'd3348;
            {7'd27,7'd125}:		p = 14'd3375;
            {7'd27,7'd126}:		p = 14'd3402;
            {7'd27,7'd127}:		p = 14'd3429;
            {7'd28,7'd0}:		p = 14'd0;
            {7'd28,7'd1}:		p = 14'd28;
            {7'd28,7'd2}:		p = 14'd56;
            {7'd28,7'd3}:		p = 14'd84;
            {7'd28,7'd4}:		p = 14'd112;
            {7'd28,7'd5}:		p = 14'd140;
            {7'd28,7'd6}:		p = 14'd168;
            {7'd28,7'd7}:		p = 14'd196;
            {7'd28,7'd8}:		p = 14'd224;
            {7'd28,7'd9}:		p = 14'd252;
            {7'd28,7'd10}:		p = 14'd280;
            {7'd28,7'd11}:		p = 14'd308;
            {7'd28,7'd12}:		p = 14'd336;
            {7'd28,7'd13}:		p = 14'd364;
            {7'd28,7'd14}:		p = 14'd392;
            {7'd28,7'd15}:		p = 14'd420;
            {7'd28,7'd16}:		p = 14'd448;
            {7'd28,7'd17}:		p = 14'd476;
            {7'd28,7'd18}:		p = 14'd504;
            {7'd28,7'd19}:		p = 14'd532;
            {7'd28,7'd20}:		p = 14'd560;
            {7'd28,7'd21}:		p = 14'd588;
            {7'd28,7'd22}:		p = 14'd616;
            {7'd28,7'd23}:		p = 14'd644;
            {7'd28,7'd24}:		p = 14'd672;
            {7'd28,7'd25}:		p = 14'd700;
            {7'd28,7'd26}:		p = 14'd728;
            {7'd28,7'd27}:		p = 14'd756;
            {7'd28,7'd28}:		p = 14'd784;
            {7'd28,7'd29}:		p = 14'd812;
            {7'd28,7'd30}:		p = 14'd840;
            {7'd28,7'd31}:		p = 14'd868;
            {7'd28,7'd32}:		p = 14'd896;
            {7'd28,7'd33}:		p = 14'd924;
            {7'd28,7'd34}:		p = 14'd952;
            {7'd28,7'd35}:		p = 14'd980;
            {7'd28,7'd36}:		p = 14'd1008;
            {7'd28,7'd37}:		p = 14'd1036;
            {7'd28,7'd38}:		p = 14'd1064;
            {7'd28,7'd39}:		p = 14'd1092;
            {7'd28,7'd40}:		p = 14'd1120;
            {7'd28,7'd41}:		p = 14'd1148;
            {7'd28,7'd42}:		p = 14'd1176;
            {7'd28,7'd43}:		p = 14'd1204;
            {7'd28,7'd44}:		p = 14'd1232;
            {7'd28,7'd45}:		p = 14'd1260;
            {7'd28,7'd46}:		p = 14'd1288;
            {7'd28,7'd47}:		p = 14'd1316;
            {7'd28,7'd48}:		p = 14'd1344;
            {7'd28,7'd49}:		p = 14'd1372;
            {7'd28,7'd50}:		p = 14'd1400;
            {7'd28,7'd51}:		p = 14'd1428;
            {7'd28,7'd52}:		p = 14'd1456;
            {7'd28,7'd53}:		p = 14'd1484;
            {7'd28,7'd54}:		p = 14'd1512;
            {7'd28,7'd55}:		p = 14'd1540;
            {7'd28,7'd56}:		p = 14'd1568;
            {7'd28,7'd57}:		p = 14'd1596;
            {7'd28,7'd58}:		p = 14'd1624;
            {7'd28,7'd59}:		p = 14'd1652;
            {7'd28,7'd60}:		p = 14'd1680;
            {7'd28,7'd61}:		p = 14'd1708;
            {7'd28,7'd62}:		p = 14'd1736;
            {7'd28,7'd63}:		p = 14'd1764;
            {7'd28,7'd64}:		p = 14'd1792;
            {7'd28,7'd65}:		p = 14'd1820;
            {7'd28,7'd66}:		p = 14'd1848;
            {7'd28,7'd67}:		p = 14'd1876;
            {7'd28,7'd68}:		p = 14'd1904;
            {7'd28,7'd69}:		p = 14'd1932;
            {7'd28,7'd70}:		p = 14'd1960;
            {7'd28,7'd71}:		p = 14'd1988;
            {7'd28,7'd72}:		p = 14'd2016;
            {7'd28,7'd73}:		p = 14'd2044;
            {7'd28,7'd74}:		p = 14'd2072;
            {7'd28,7'd75}:		p = 14'd2100;
            {7'd28,7'd76}:		p = 14'd2128;
            {7'd28,7'd77}:		p = 14'd2156;
            {7'd28,7'd78}:		p = 14'd2184;
            {7'd28,7'd79}:		p = 14'd2212;
            {7'd28,7'd80}:		p = 14'd2240;
            {7'd28,7'd81}:		p = 14'd2268;
            {7'd28,7'd82}:		p = 14'd2296;
            {7'd28,7'd83}:		p = 14'd2324;
            {7'd28,7'd84}:		p = 14'd2352;
            {7'd28,7'd85}:		p = 14'd2380;
            {7'd28,7'd86}:		p = 14'd2408;
            {7'd28,7'd87}:		p = 14'd2436;
            {7'd28,7'd88}:		p = 14'd2464;
            {7'd28,7'd89}:		p = 14'd2492;
            {7'd28,7'd90}:		p = 14'd2520;
            {7'd28,7'd91}:		p = 14'd2548;
            {7'd28,7'd92}:		p = 14'd2576;
            {7'd28,7'd93}:		p = 14'd2604;
            {7'd28,7'd94}:		p = 14'd2632;
            {7'd28,7'd95}:		p = 14'd2660;
            {7'd28,7'd96}:		p = 14'd2688;
            {7'd28,7'd97}:		p = 14'd2716;
            {7'd28,7'd98}:		p = 14'd2744;
            {7'd28,7'd99}:		p = 14'd2772;
            {7'd28,7'd100}:		p = 14'd2800;
            {7'd28,7'd101}:		p = 14'd2828;
            {7'd28,7'd102}:		p = 14'd2856;
            {7'd28,7'd103}:		p = 14'd2884;
            {7'd28,7'd104}:		p = 14'd2912;
            {7'd28,7'd105}:		p = 14'd2940;
            {7'd28,7'd106}:		p = 14'd2968;
            {7'd28,7'd107}:		p = 14'd2996;
            {7'd28,7'd108}:		p = 14'd3024;
            {7'd28,7'd109}:		p = 14'd3052;
            {7'd28,7'd110}:		p = 14'd3080;
            {7'd28,7'd111}:		p = 14'd3108;
            {7'd28,7'd112}:		p = 14'd3136;
            {7'd28,7'd113}:		p = 14'd3164;
            {7'd28,7'd114}:		p = 14'd3192;
            {7'd28,7'd115}:		p = 14'd3220;
            {7'd28,7'd116}:		p = 14'd3248;
            {7'd28,7'd117}:		p = 14'd3276;
            {7'd28,7'd118}:		p = 14'd3304;
            {7'd28,7'd119}:		p = 14'd3332;
            {7'd28,7'd120}:		p = 14'd3360;
            {7'd28,7'd121}:		p = 14'd3388;
            {7'd28,7'd122}:		p = 14'd3416;
            {7'd28,7'd123}:		p = 14'd3444;
            {7'd28,7'd124}:		p = 14'd3472;
            {7'd28,7'd125}:		p = 14'd3500;
            {7'd28,7'd126}:		p = 14'd3528;
            {7'd28,7'd127}:		p = 14'd3556;
            {7'd29,7'd0}:		p = 14'd0;
            {7'd29,7'd1}:		p = 14'd29;
            {7'd29,7'd2}:		p = 14'd58;
            {7'd29,7'd3}:		p = 14'd87;
            {7'd29,7'd4}:		p = 14'd116;
            {7'd29,7'd5}:		p = 14'd145;
            {7'd29,7'd6}:		p = 14'd174;
            {7'd29,7'd7}:		p = 14'd203;
            {7'd29,7'd8}:		p = 14'd232;
            {7'd29,7'd9}:		p = 14'd261;
            {7'd29,7'd10}:		p = 14'd290;
            {7'd29,7'd11}:		p = 14'd319;
            {7'd29,7'd12}:		p = 14'd348;
            {7'd29,7'd13}:		p = 14'd377;
            {7'd29,7'd14}:		p = 14'd406;
            {7'd29,7'd15}:		p = 14'd435;
            {7'd29,7'd16}:		p = 14'd464;
            {7'd29,7'd17}:		p = 14'd493;
            {7'd29,7'd18}:		p = 14'd522;
            {7'd29,7'd19}:		p = 14'd551;
            {7'd29,7'd20}:		p = 14'd580;
            {7'd29,7'd21}:		p = 14'd609;
            {7'd29,7'd22}:		p = 14'd638;
            {7'd29,7'd23}:		p = 14'd667;
            {7'd29,7'd24}:		p = 14'd696;
            {7'd29,7'd25}:		p = 14'd725;
            {7'd29,7'd26}:		p = 14'd754;
            {7'd29,7'd27}:		p = 14'd783;
            {7'd29,7'd28}:		p = 14'd812;
            {7'd29,7'd29}:		p = 14'd841;
            {7'd29,7'd30}:		p = 14'd870;
            {7'd29,7'd31}:		p = 14'd899;
            {7'd29,7'd32}:		p = 14'd928;
            {7'd29,7'd33}:		p = 14'd957;
            {7'd29,7'd34}:		p = 14'd986;
            {7'd29,7'd35}:		p = 14'd1015;
            {7'd29,7'd36}:		p = 14'd1044;
            {7'd29,7'd37}:		p = 14'd1073;
            {7'd29,7'd38}:		p = 14'd1102;
            {7'd29,7'd39}:		p = 14'd1131;
            {7'd29,7'd40}:		p = 14'd1160;
            {7'd29,7'd41}:		p = 14'd1189;
            {7'd29,7'd42}:		p = 14'd1218;
            {7'd29,7'd43}:		p = 14'd1247;
            {7'd29,7'd44}:		p = 14'd1276;
            {7'd29,7'd45}:		p = 14'd1305;
            {7'd29,7'd46}:		p = 14'd1334;
            {7'd29,7'd47}:		p = 14'd1363;
            {7'd29,7'd48}:		p = 14'd1392;
            {7'd29,7'd49}:		p = 14'd1421;
            {7'd29,7'd50}:		p = 14'd1450;
            {7'd29,7'd51}:		p = 14'd1479;
            {7'd29,7'd52}:		p = 14'd1508;
            {7'd29,7'd53}:		p = 14'd1537;
            {7'd29,7'd54}:		p = 14'd1566;
            {7'd29,7'd55}:		p = 14'd1595;
            {7'd29,7'd56}:		p = 14'd1624;
            {7'd29,7'd57}:		p = 14'd1653;
            {7'd29,7'd58}:		p = 14'd1682;
            {7'd29,7'd59}:		p = 14'd1711;
            {7'd29,7'd60}:		p = 14'd1740;
            {7'd29,7'd61}:		p = 14'd1769;
            {7'd29,7'd62}:		p = 14'd1798;
            {7'd29,7'd63}:		p = 14'd1827;
            {7'd29,7'd64}:		p = 14'd1856;
            {7'd29,7'd65}:		p = 14'd1885;
            {7'd29,7'd66}:		p = 14'd1914;
            {7'd29,7'd67}:		p = 14'd1943;
            {7'd29,7'd68}:		p = 14'd1972;
            {7'd29,7'd69}:		p = 14'd2001;
            {7'd29,7'd70}:		p = 14'd2030;
            {7'd29,7'd71}:		p = 14'd2059;
            {7'd29,7'd72}:		p = 14'd2088;
            {7'd29,7'd73}:		p = 14'd2117;
            {7'd29,7'd74}:		p = 14'd2146;
            {7'd29,7'd75}:		p = 14'd2175;
            {7'd29,7'd76}:		p = 14'd2204;
            {7'd29,7'd77}:		p = 14'd2233;
            {7'd29,7'd78}:		p = 14'd2262;
            {7'd29,7'd79}:		p = 14'd2291;
            {7'd29,7'd80}:		p = 14'd2320;
            {7'd29,7'd81}:		p = 14'd2349;
            {7'd29,7'd82}:		p = 14'd2378;
            {7'd29,7'd83}:		p = 14'd2407;
            {7'd29,7'd84}:		p = 14'd2436;
            {7'd29,7'd85}:		p = 14'd2465;
            {7'd29,7'd86}:		p = 14'd2494;
            {7'd29,7'd87}:		p = 14'd2523;
            {7'd29,7'd88}:		p = 14'd2552;
            {7'd29,7'd89}:		p = 14'd2581;
            {7'd29,7'd90}:		p = 14'd2610;
            {7'd29,7'd91}:		p = 14'd2639;
            {7'd29,7'd92}:		p = 14'd2668;
            {7'd29,7'd93}:		p = 14'd2697;
            {7'd29,7'd94}:		p = 14'd2726;
            {7'd29,7'd95}:		p = 14'd2755;
            {7'd29,7'd96}:		p = 14'd2784;
            {7'd29,7'd97}:		p = 14'd2813;
            {7'd29,7'd98}:		p = 14'd2842;
            {7'd29,7'd99}:		p = 14'd2871;
            {7'd29,7'd100}:		p = 14'd2900;
            {7'd29,7'd101}:		p = 14'd2929;
            {7'd29,7'd102}:		p = 14'd2958;
            {7'd29,7'd103}:		p = 14'd2987;
            {7'd29,7'd104}:		p = 14'd3016;
            {7'd29,7'd105}:		p = 14'd3045;
            {7'd29,7'd106}:		p = 14'd3074;
            {7'd29,7'd107}:		p = 14'd3103;
            {7'd29,7'd108}:		p = 14'd3132;
            {7'd29,7'd109}:		p = 14'd3161;
            {7'd29,7'd110}:		p = 14'd3190;
            {7'd29,7'd111}:		p = 14'd3219;
            {7'd29,7'd112}:		p = 14'd3248;
            {7'd29,7'd113}:		p = 14'd3277;
            {7'd29,7'd114}:		p = 14'd3306;
            {7'd29,7'd115}:		p = 14'd3335;
            {7'd29,7'd116}:		p = 14'd3364;
            {7'd29,7'd117}:		p = 14'd3393;
            {7'd29,7'd118}:		p = 14'd3422;
            {7'd29,7'd119}:		p = 14'd3451;
            {7'd29,7'd120}:		p = 14'd3480;
            {7'd29,7'd121}:		p = 14'd3509;
            {7'd29,7'd122}:		p = 14'd3538;
            {7'd29,7'd123}:		p = 14'd3567;
            {7'd29,7'd124}:		p = 14'd3596;
            {7'd29,7'd125}:		p = 14'd3625;
            {7'd29,7'd126}:		p = 14'd3654;
            {7'd29,7'd127}:		p = 14'd3683;
            {7'd30,7'd0}:		p = 14'd0;
            {7'd30,7'd1}:		p = 14'd30;
            {7'd30,7'd2}:		p = 14'd60;
            {7'd30,7'd3}:		p = 14'd90;
            {7'd30,7'd4}:		p = 14'd120;
            {7'd30,7'd5}:		p = 14'd150;
            {7'd30,7'd6}:		p = 14'd180;
            {7'd30,7'd7}:		p = 14'd210;
            {7'd30,7'd8}:		p = 14'd240;
            {7'd30,7'd9}:		p = 14'd270;
            {7'd30,7'd10}:		p = 14'd300;
            {7'd30,7'd11}:		p = 14'd330;
            {7'd30,7'd12}:		p = 14'd360;
            {7'd30,7'd13}:		p = 14'd390;
            {7'd30,7'd14}:		p = 14'd420;
            {7'd30,7'd15}:		p = 14'd450;
            {7'd30,7'd16}:		p = 14'd480;
            {7'd30,7'd17}:		p = 14'd510;
            {7'd30,7'd18}:		p = 14'd540;
            {7'd30,7'd19}:		p = 14'd570;
            {7'd30,7'd20}:		p = 14'd600;
            {7'd30,7'd21}:		p = 14'd630;
            {7'd30,7'd22}:		p = 14'd660;
            {7'd30,7'd23}:		p = 14'd690;
            {7'd30,7'd24}:		p = 14'd720;
            {7'd30,7'd25}:		p = 14'd750;
            {7'd30,7'd26}:		p = 14'd780;
            {7'd30,7'd27}:		p = 14'd810;
            {7'd30,7'd28}:		p = 14'd840;
            {7'd30,7'd29}:		p = 14'd870;
            {7'd30,7'd30}:		p = 14'd900;
            {7'd30,7'd31}:		p = 14'd930;
            {7'd30,7'd32}:		p = 14'd960;
            {7'd30,7'd33}:		p = 14'd990;
            {7'd30,7'd34}:		p = 14'd1020;
            {7'd30,7'd35}:		p = 14'd1050;
            {7'd30,7'd36}:		p = 14'd1080;
            {7'd30,7'd37}:		p = 14'd1110;
            {7'd30,7'd38}:		p = 14'd1140;
            {7'd30,7'd39}:		p = 14'd1170;
            {7'd30,7'd40}:		p = 14'd1200;
            {7'd30,7'd41}:		p = 14'd1230;
            {7'd30,7'd42}:		p = 14'd1260;
            {7'd30,7'd43}:		p = 14'd1290;
            {7'd30,7'd44}:		p = 14'd1320;
            {7'd30,7'd45}:		p = 14'd1350;
            {7'd30,7'd46}:		p = 14'd1380;
            {7'd30,7'd47}:		p = 14'd1410;
            {7'd30,7'd48}:		p = 14'd1440;
            {7'd30,7'd49}:		p = 14'd1470;
            {7'd30,7'd50}:		p = 14'd1500;
            {7'd30,7'd51}:		p = 14'd1530;
            {7'd30,7'd52}:		p = 14'd1560;
            {7'd30,7'd53}:		p = 14'd1590;
            {7'd30,7'd54}:		p = 14'd1620;
            {7'd30,7'd55}:		p = 14'd1650;
            {7'd30,7'd56}:		p = 14'd1680;
            {7'd30,7'd57}:		p = 14'd1710;
            {7'd30,7'd58}:		p = 14'd1740;
            {7'd30,7'd59}:		p = 14'd1770;
            {7'd30,7'd60}:		p = 14'd1800;
            {7'd30,7'd61}:		p = 14'd1830;
            {7'd30,7'd62}:		p = 14'd1860;
            {7'd30,7'd63}:		p = 14'd1890;
            {7'd30,7'd64}:		p = 14'd1920;
            {7'd30,7'd65}:		p = 14'd1950;
            {7'd30,7'd66}:		p = 14'd1980;
            {7'd30,7'd67}:		p = 14'd2010;
            {7'd30,7'd68}:		p = 14'd2040;
            {7'd30,7'd69}:		p = 14'd2070;
            {7'd30,7'd70}:		p = 14'd2100;
            {7'd30,7'd71}:		p = 14'd2130;
            {7'd30,7'd72}:		p = 14'd2160;
            {7'd30,7'd73}:		p = 14'd2190;
            {7'd30,7'd74}:		p = 14'd2220;
            {7'd30,7'd75}:		p = 14'd2250;
            {7'd30,7'd76}:		p = 14'd2280;
            {7'd30,7'd77}:		p = 14'd2310;
            {7'd30,7'd78}:		p = 14'd2340;
            {7'd30,7'd79}:		p = 14'd2370;
            {7'd30,7'd80}:		p = 14'd2400;
            {7'd30,7'd81}:		p = 14'd2430;
            {7'd30,7'd82}:		p = 14'd2460;
            {7'd30,7'd83}:		p = 14'd2490;
            {7'd30,7'd84}:		p = 14'd2520;
            {7'd30,7'd85}:		p = 14'd2550;
            {7'd30,7'd86}:		p = 14'd2580;
            {7'd30,7'd87}:		p = 14'd2610;
            {7'd30,7'd88}:		p = 14'd2640;
            {7'd30,7'd89}:		p = 14'd2670;
            {7'd30,7'd90}:		p = 14'd2700;
            {7'd30,7'd91}:		p = 14'd2730;
            {7'd30,7'd92}:		p = 14'd2760;
            {7'd30,7'd93}:		p = 14'd2790;
            {7'd30,7'd94}:		p = 14'd2820;
            {7'd30,7'd95}:		p = 14'd2850;
            {7'd30,7'd96}:		p = 14'd2880;
            {7'd30,7'd97}:		p = 14'd2910;
            {7'd30,7'd98}:		p = 14'd2940;
            {7'd30,7'd99}:		p = 14'd2970;
            {7'd30,7'd100}:		p = 14'd3000;
            {7'd30,7'd101}:		p = 14'd3030;
            {7'd30,7'd102}:		p = 14'd3060;
            {7'd30,7'd103}:		p = 14'd3090;
            {7'd30,7'd104}:		p = 14'd3120;
            {7'd30,7'd105}:		p = 14'd3150;
            {7'd30,7'd106}:		p = 14'd3180;
            {7'd30,7'd107}:		p = 14'd3210;
            {7'd30,7'd108}:		p = 14'd3240;
            {7'd30,7'd109}:		p = 14'd3270;
            {7'd30,7'd110}:		p = 14'd3300;
            {7'd30,7'd111}:		p = 14'd3330;
            {7'd30,7'd112}:		p = 14'd3360;
            {7'd30,7'd113}:		p = 14'd3390;
            {7'd30,7'd114}:		p = 14'd3420;
            {7'd30,7'd115}:		p = 14'd3450;
            {7'd30,7'd116}:		p = 14'd3480;
            {7'd30,7'd117}:		p = 14'd3510;
            {7'd30,7'd118}:		p = 14'd3540;
            {7'd30,7'd119}:		p = 14'd3570;
            {7'd30,7'd120}:		p = 14'd3600;
            {7'd30,7'd121}:		p = 14'd3630;
            {7'd30,7'd122}:		p = 14'd3660;
            {7'd30,7'd123}:		p = 14'd3690;
            {7'd30,7'd124}:		p = 14'd3720;
            {7'd30,7'd125}:		p = 14'd3750;
            {7'd30,7'd126}:		p = 14'd3780;
            {7'd30,7'd127}:		p = 14'd3810;
            {7'd31,7'd0}:		p = 14'd0;
            {7'd31,7'd1}:		p = 14'd31;
            {7'd31,7'd2}:		p = 14'd62;
            {7'd31,7'd3}:		p = 14'd93;
            {7'd31,7'd4}:		p = 14'd124;
            {7'd31,7'd5}:		p = 14'd155;
            {7'd31,7'd6}:		p = 14'd186;
            {7'd31,7'd7}:		p = 14'd217;
            {7'd31,7'd8}:		p = 14'd248;
            {7'd31,7'd9}:		p = 14'd279;
            {7'd31,7'd10}:		p = 14'd310;
            {7'd31,7'd11}:		p = 14'd341;
            {7'd31,7'd12}:		p = 14'd372;
            {7'd31,7'd13}:		p = 14'd403;
            {7'd31,7'd14}:		p = 14'd434;
            {7'd31,7'd15}:		p = 14'd465;
            {7'd31,7'd16}:		p = 14'd496;
            {7'd31,7'd17}:		p = 14'd527;
            {7'd31,7'd18}:		p = 14'd558;
            {7'd31,7'd19}:		p = 14'd589;
            {7'd31,7'd20}:		p = 14'd620;
            {7'd31,7'd21}:		p = 14'd651;
            {7'd31,7'd22}:		p = 14'd682;
            {7'd31,7'd23}:		p = 14'd713;
            {7'd31,7'd24}:		p = 14'd744;
            {7'd31,7'd25}:		p = 14'd775;
            {7'd31,7'd26}:		p = 14'd806;
            {7'd31,7'd27}:		p = 14'd837;
            {7'd31,7'd28}:		p = 14'd868;
            {7'd31,7'd29}:		p = 14'd899;
            {7'd31,7'd30}:		p = 14'd930;
            {7'd31,7'd31}:		p = 14'd961;
            {7'd31,7'd32}:		p = 14'd992;
            {7'd31,7'd33}:		p = 14'd1023;
            {7'd31,7'd34}:		p = 14'd1054;
            {7'd31,7'd35}:		p = 14'd1085;
            {7'd31,7'd36}:		p = 14'd1116;
            {7'd31,7'd37}:		p = 14'd1147;
            {7'd31,7'd38}:		p = 14'd1178;
            {7'd31,7'd39}:		p = 14'd1209;
            {7'd31,7'd40}:		p = 14'd1240;
            {7'd31,7'd41}:		p = 14'd1271;
            {7'd31,7'd42}:		p = 14'd1302;
            {7'd31,7'd43}:		p = 14'd1333;
            {7'd31,7'd44}:		p = 14'd1364;
            {7'd31,7'd45}:		p = 14'd1395;
            {7'd31,7'd46}:		p = 14'd1426;
            {7'd31,7'd47}:		p = 14'd1457;
            {7'd31,7'd48}:		p = 14'd1488;
            {7'd31,7'd49}:		p = 14'd1519;
            {7'd31,7'd50}:		p = 14'd1550;
            {7'd31,7'd51}:		p = 14'd1581;
            {7'd31,7'd52}:		p = 14'd1612;
            {7'd31,7'd53}:		p = 14'd1643;
            {7'd31,7'd54}:		p = 14'd1674;
            {7'd31,7'd55}:		p = 14'd1705;
            {7'd31,7'd56}:		p = 14'd1736;
            {7'd31,7'd57}:		p = 14'd1767;
            {7'd31,7'd58}:		p = 14'd1798;
            {7'd31,7'd59}:		p = 14'd1829;
            {7'd31,7'd60}:		p = 14'd1860;
            {7'd31,7'd61}:		p = 14'd1891;
            {7'd31,7'd62}:		p = 14'd1922;
            {7'd31,7'd63}:		p = 14'd1953;
            {7'd31,7'd64}:		p = 14'd1984;
            {7'd31,7'd65}:		p = 14'd2015;
            {7'd31,7'd66}:		p = 14'd2046;
            {7'd31,7'd67}:		p = 14'd2077;
            {7'd31,7'd68}:		p = 14'd2108;
            {7'd31,7'd69}:		p = 14'd2139;
            {7'd31,7'd70}:		p = 14'd2170;
            {7'd31,7'd71}:		p = 14'd2201;
            {7'd31,7'd72}:		p = 14'd2232;
            {7'd31,7'd73}:		p = 14'd2263;
            {7'd31,7'd74}:		p = 14'd2294;
            {7'd31,7'd75}:		p = 14'd2325;
            {7'd31,7'd76}:		p = 14'd2356;
            {7'd31,7'd77}:		p = 14'd2387;
            {7'd31,7'd78}:		p = 14'd2418;
            {7'd31,7'd79}:		p = 14'd2449;
            {7'd31,7'd80}:		p = 14'd2480;
            {7'd31,7'd81}:		p = 14'd2511;
            {7'd31,7'd82}:		p = 14'd2542;
            {7'd31,7'd83}:		p = 14'd2573;
            {7'd31,7'd84}:		p = 14'd2604;
            {7'd31,7'd85}:		p = 14'd2635;
            {7'd31,7'd86}:		p = 14'd2666;
            {7'd31,7'd87}:		p = 14'd2697;
            {7'd31,7'd88}:		p = 14'd2728;
            {7'd31,7'd89}:		p = 14'd2759;
            {7'd31,7'd90}:		p = 14'd2790;
            {7'd31,7'd91}:		p = 14'd2821;
            {7'd31,7'd92}:		p = 14'd2852;
            {7'd31,7'd93}:		p = 14'd2883;
            {7'd31,7'd94}:		p = 14'd2914;
            {7'd31,7'd95}:		p = 14'd2945;
            {7'd31,7'd96}:		p = 14'd2976;
            {7'd31,7'd97}:		p = 14'd3007;
            {7'd31,7'd98}:		p = 14'd3038;
            {7'd31,7'd99}:		p = 14'd3069;
            {7'd31,7'd100}:		p = 14'd3100;
            {7'd31,7'd101}:		p = 14'd3131;
            {7'd31,7'd102}:		p = 14'd3162;
            {7'd31,7'd103}:		p = 14'd3193;
            {7'd31,7'd104}:		p = 14'd3224;
            {7'd31,7'd105}:		p = 14'd3255;
            {7'd31,7'd106}:		p = 14'd3286;
            {7'd31,7'd107}:		p = 14'd3317;
            {7'd31,7'd108}:		p = 14'd3348;
            {7'd31,7'd109}:		p = 14'd3379;
            {7'd31,7'd110}:		p = 14'd3410;
            {7'd31,7'd111}:		p = 14'd3441;
            {7'd31,7'd112}:		p = 14'd3472;
            {7'd31,7'd113}:		p = 14'd3503;
            {7'd31,7'd114}:		p = 14'd3534;
            {7'd31,7'd115}:		p = 14'd3565;
            {7'd31,7'd116}:		p = 14'd3596;
            {7'd31,7'd117}:		p = 14'd3627;
            {7'd31,7'd118}:		p = 14'd3658;
            {7'd31,7'd119}:		p = 14'd3689;
            {7'd31,7'd120}:		p = 14'd3720;
            {7'd31,7'd121}:		p = 14'd3751;
            {7'd31,7'd122}:		p = 14'd3782;
            {7'd31,7'd123}:		p = 14'd3813;
            {7'd31,7'd124}:		p = 14'd3844;
            {7'd31,7'd125}:		p = 14'd3875;
            {7'd31,7'd126}:		p = 14'd3906;
            {7'd31,7'd127}:		p = 14'd3937;
            {7'd32,7'd0}:		p = 14'd0;
            {7'd32,7'd1}:		p = 14'd32;
            {7'd32,7'd2}:		p = 14'd64;
            {7'd32,7'd3}:		p = 14'd96;
            {7'd32,7'd4}:		p = 14'd128;
            {7'd32,7'd5}:		p = 14'd160;
            {7'd32,7'd6}:		p = 14'd192;
            {7'd32,7'd7}:		p = 14'd224;
            {7'd32,7'd8}:		p = 14'd256;
            {7'd32,7'd9}:		p = 14'd288;
            {7'd32,7'd10}:		p = 14'd320;
            {7'd32,7'd11}:		p = 14'd352;
            {7'd32,7'd12}:		p = 14'd384;
            {7'd32,7'd13}:		p = 14'd416;
            {7'd32,7'd14}:		p = 14'd448;
            {7'd32,7'd15}:		p = 14'd480;
            {7'd32,7'd16}:		p = 14'd512;
            {7'd32,7'd17}:		p = 14'd544;
            {7'd32,7'd18}:		p = 14'd576;
            {7'd32,7'd19}:		p = 14'd608;
            {7'd32,7'd20}:		p = 14'd640;
            {7'd32,7'd21}:		p = 14'd672;
            {7'd32,7'd22}:		p = 14'd704;
            {7'd32,7'd23}:		p = 14'd736;
            {7'd32,7'd24}:		p = 14'd768;
            {7'd32,7'd25}:		p = 14'd800;
            {7'd32,7'd26}:		p = 14'd832;
            {7'd32,7'd27}:		p = 14'd864;
            {7'd32,7'd28}:		p = 14'd896;
            {7'd32,7'd29}:		p = 14'd928;
            {7'd32,7'd30}:		p = 14'd960;
            {7'd32,7'd31}:		p = 14'd992;
            {7'd32,7'd32}:		p = 14'd1024;
            {7'd32,7'd33}:		p = 14'd1056;
            {7'd32,7'd34}:		p = 14'd1088;
            {7'd32,7'd35}:		p = 14'd1120;
            {7'd32,7'd36}:		p = 14'd1152;
            {7'd32,7'd37}:		p = 14'd1184;
            {7'd32,7'd38}:		p = 14'd1216;
            {7'd32,7'd39}:		p = 14'd1248;
            {7'd32,7'd40}:		p = 14'd1280;
            {7'd32,7'd41}:		p = 14'd1312;
            {7'd32,7'd42}:		p = 14'd1344;
            {7'd32,7'd43}:		p = 14'd1376;
            {7'd32,7'd44}:		p = 14'd1408;
            {7'd32,7'd45}:		p = 14'd1440;
            {7'd32,7'd46}:		p = 14'd1472;
            {7'd32,7'd47}:		p = 14'd1504;
            {7'd32,7'd48}:		p = 14'd1536;
            {7'd32,7'd49}:		p = 14'd1568;
            {7'd32,7'd50}:		p = 14'd1600;
            {7'd32,7'd51}:		p = 14'd1632;
            {7'd32,7'd52}:		p = 14'd1664;
            {7'd32,7'd53}:		p = 14'd1696;
            {7'd32,7'd54}:		p = 14'd1728;
            {7'd32,7'd55}:		p = 14'd1760;
            {7'd32,7'd56}:		p = 14'd1792;
            {7'd32,7'd57}:		p = 14'd1824;
            {7'd32,7'd58}:		p = 14'd1856;
            {7'd32,7'd59}:		p = 14'd1888;
            {7'd32,7'd60}:		p = 14'd1920;
            {7'd32,7'd61}:		p = 14'd1952;
            {7'd32,7'd62}:		p = 14'd1984;
            {7'd32,7'd63}:		p = 14'd2016;
            {7'd32,7'd64}:		p = 14'd2048;
            {7'd32,7'd65}:		p = 14'd2080;
            {7'd32,7'd66}:		p = 14'd2112;
            {7'd32,7'd67}:		p = 14'd2144;
            {7'd32,7'd68}:		p = 14'd2176;
            {7'd32,7'd69}:		p = 14'd2208;
            {7'd32,7'd70}:		p = 14'd2240;
            {7'd32,7'd71}:		p = 14'd2272;
            {7'd32,7'd72}:		p = 14'd2304;
            {7'd32,7'd73}:		p = 14'd2336;
            {7'd32,7'd74}:		p = 14'd2368;
            {7'd32,7'd75}:		p = 14'd2400;
            {7'd32,7'd76}:		p = 14'd2432;
            {7'd32,7'd77}:		p = 14'd2464;
            {7'd32,7'd78}:		p = 14'd2496;
            {7'd32,7'd79}:		p = 14'd2528;
            {7'd32,7'd80}:		p = 14'd2560;
            {7'd32,7'd81}:		p = 14'd2592;
            {7'd32,7'd82}:		p = 14'd2624;
            {7'd32,7'd83}:		p = 14'd2656;
            {7'd32,7'd84}:		p = 14'd2688;
            {7'd32,7'd85}:		p = 14'd2720;
            {7'd32,7'd86}:		p = 14'd2752;
            {7'd32,7'd87}:		p = 14'd2784;
            {7'd32,7'd88}:		p = 14'd2816;
            {7'd32,7'd89}:		p = 14'd2848;
            {7'd32,7'd90}:		p = 14'd2880;
            {7'd32,7'd91}:		p = 14'd2912;
            {7'd32,7'd92}:		p = 14'd2944;
            {7'd32,7'd93}:		p = 14'd2976;
            {7'd32,7'd94}:		p = 14'd3008;
            {7'd32,7'd95}:		p = 14'd3040;
            {7'd32,7'd96}:		p = 14'd3072;
            {7'd32,7'd97}:		p = 14'd3104;
            {7'd32,7'd98}:		p = 14'd3136;
            {7'd32,7'd99}:		p = 14'd3168;
            {7'd32,7'd100}:		p = 14'd3200;
            {7'd32,7'd101}:		p = 14'd3232;
            {7'd32,7'd102}:		p = 14'd3264;
            {7'd32,7'd103}:		p = 14'd3296;
            {7'd32,7'd104}:		p = 14'd3328;
            {7'd32,7'd105}:		p = 14'd3360;
            {7'd32,7'd106}:		p = 14'd3392;
            {7'd32,7'd107}:		p = 14'd3424;
            {7'd32,7'd108}:		p = 14'd3456;
            {7'd32,7'd109}:		p = 14'd3488;
            {7'd32,7'd110}:		p = 14'd3520;
            {7'd32,7'd111}:		p = 14'd3552;
            {7'd32,7'd112}:		p = 14'd3584;
            {7'd32,7'd113}:		p = 14'd3616;
            {7'd32,7'd114}:		p = 14'd3648;
            {7'd32,7'd115}:		p = 14'd3680;
            {7'd32,7'd116}:		p = 14'd3712;
            {7'd32,7'd117}:		p = 14'd3744;
            {7'd32,7'd118}:		p = 14'd3776;
            {7'd32,7'd119}:		p = 14'd3808;
            {7'd32,7'd120}:		p = 14'd3840;
            {7'd32,7'd121}:		p = 14'd3872;
            {7'd32,7'd122}:		p = 14'd3904;
            {7'd32,7'd123}:		p = 14'd3936;
            {7'd32,7'd124}:		p = 14'd3968;
            {7'd32,7'd125}:		p = 14'd4000;
            {7'd32,7'd126}:		p = 14'd4032;
            {7'd32,7'd127}:		p = 14'd4064;
            {7'd33,7'd0}:		p = 14'd0;
            {7'd33,7'd1}:		p = 14'd33;
            {7'd33,7'd2}:		p = 14'd66;
            {7'd33,7'd3}:		p = 14'd99;
            {7'd33,7'd4}:		p = 14'd132;
            {7'd33,7'd5}:		p = 14'd165;
            {7'd33,7'd6}:		p = 14'd198;
            {7'd33,7'd7}:		p = 14'd231;
            {7'd33,7'd8}:		p = 14'd264;
            {7'd33,7'd9}:		p = 14'd297;
            {7'd33,7'd10}:		p = 14'd330;
            {7'd33,7'd11}:		p = 14'd363;
            {7'd33,7'd12}:		p = 14'd396;
            {7'd33,7'd13}:		p = 14'd429;
            {7'd33,7'd14}:		p = 14'd462;
            {7'd33,7'd15}:		p = 14'd495;
            {7'd33,7'd16}:		p = 14'd528;
            {7'd33,7'd17}:		p = 14'd561;
            {7'd33,7'd18}:		p = 14'd594;
            {7'd33,7'd19}:		p = 14'd627;
            {7'd33,7'd20}:		p = 14'd660;
            {7'd33,7'd21}:		p = 14'd693;
            {7'd33,7'd22}:		p = 14'd726;
            {7'd33,7'd23}:		p = 14'd759;
            {7'd33,7'd24}:		p = 14'd792;
            {7'd33,7'd25}:		p = 14'd825;
            {7'd33,7'd26}:		p = 14'd858;
            {7'd33,7'd27}:		p = 14'd891;
            {7'd33,7'd28}:		p = 14'd924;
            {7'd33,7'd29}:		p = 14'd957;
            {7'd33,7'd30}:		p = 14'd990;
            {7'd33,7'd31}:		p = 14'd1023;
            {7'd33,7'd32}:		p = 14'd1056;
            {7'd33,7'd33}:		p = 14'd1089;
            {7'd33,7'd34}:		p = 14'd1122;
            {7'd33,7'd35}:		p = 14'd1155;
            {7'd33,7'd36}:		p = 14'd1188;
            {7'd33,7'd37}:		p = 14'd1221;
            {7'd33,7'd38}:		p = 14'd1254;
            {7'd33,7'd39}:		p = 14'd1287;
            {7'd33,7'd40}:		p = 14'd1320;
            {7'd33,7'd41}:		p = 14'd1353;
            {7'd33,7'd42}:		p = 14'd1386;
            {7'd33,7'd43}:		p = 14'd1419;
            {7'd33,7'd44}:		p = 14'd1452;
            {7'd33,7'd45}:		p = 14'd1485;
            {7'd33,7'd46}:		p = 14'd1518;
            {7'd33,7'd47}:		p = 14'd1551;
            {7'd33,7'd48}:		p = 14'd1584;
            {7'd33,7'd49}:		p = 14'd1617;
            {7'd33,7'd50}:		p = 14'd1650;
            {7'd33,7'd51}:		p = 14'd1683;
            {7'd33,7'd52}:		p = 14'd1716;
            {7'd33,7'd53}:		p = 14'd1749;
            {7'd33,7'd54}:		p = 14'd1782;
            {7'd33,7'd55}:		p = 14'd1815;
            {7'd33,7'd56}:		p = 14'd1848;
            {7'd33,7'd57}:		p = 14'd1881;
            {7'd33,7'd58}:		p = 14'd1914;
            {7'd33,7'd59}:		p = 14'd1947;
            {7'd33,7'd60}:		p = 14'd1980;
            {7'd33,7'd61}:		p = 14'd2013;
            {7'd33,7'd62}:		p = 14'd2046;
            {7'd33,7'd63}:		p = 14'd2079;
            {7'd33,7'd64}:		p = 14'd2112;
            {7'd33,7'd65}:		p = 14'd2145;
            {7'd33,7'd66}:		p = 14'd2178;
            {7'd33,7'd67}:		p = 14'd2211;
            {7'd33,7'd68}:		p = 14'd2244;
            {7'd33,7'd69}:		p = 14'd2277;
            {7'd33,7'd70}:		p = 14'd2310;
            {7'd33,7'd71}:		p = 14'd2343;
            {7'd33,7'd72}:		p = 14'd2376;
            {7'd33,7'd73}:		p = 14'd2409;
            {7'd33,7'd74}:		p = 14'd2442;
            {7'd33,7'd75}:		p = 14'd2475;
            {7'd33,7'd76}:		p = 14'd2508;
            {7'd33,7'd77}:		p = 14'd2541;
            {7'd33,7'd78}:		p = 14'd2574;
            {7'd33,7'd79}:		p = 14'd2607;
            {7'd33,7'd80}:		p = 14'd2640;
            {7'd33,7'd81}:		p = 14'd2673;
            {7'd33,7'd82}:		p = 14'd2706;
            {7'd33,7'd83}:		p = 14'd2739;
            {7'd33,7'd84}:		p = 14'd2772;
            {7'd33,7'd85}:		p = 14'd2805;
            {7'd33,7'd86}:		p = 14'd2838;
            {7'd33,7'd87}:		p = 14'd2871;
            {7'd33,7'd88}:		p = 14'd2904;
            {7'd33,7'd89}:		p = 14'd2937;
            {7'd33,7'd90}:		p = 14'd2970;
            {7'd33,7'd91}:		p = 14'd3003;
            {7'd33,7'd92}:		p = 14'd3036;
            {7'd33,7'd93}:		p = 14'd3069;
            {7'd33,7'd94}:		p = 14'd3102;
            {7'd33,7'd95}:		p = 14'd3135;
            {7'd33,7'd96}:		p = 14'd3168;
            {7'd33,7'd97}:		p = 14'd3201;
            {7'd33,7'd98}:		p = 14'd3234;
            {7'd33,7'd99}:		p = 14'd3267;
            {7'd33,7'd100}:		p = 14'd3300;
            {7'd33,7'd101}:		p = 14'd3333;
            {7'd33,7'd102}:		p = 14'd3366;
            {7'd33,7'd103}:		p = 14'd3399;
            {7'd33,7'd104}:		p = 14'd3432;
            {7'd33,7'd105}:		p = 14'd3465;
            {7'd33,7'd106}:		p = 14'd3498;
            {7'd33,7'd107}:		p = 14'd3531;
            {7'd33,7'd108}:		p = 14'd3564;
            {7'd33,7'd109}:		p = 14'd3597;
            {7'd33,7'd110}:		p = 14'd3630;
            {7'd33,7'd111}:		p = 14'd3663;
            {7'd33,7'd112}:		p = 14'd3696;
            {7'd33,7'd113}:		p = 14'd3729;
            {7'd33,7'd114}:		p = 14'd3762;
            {7'd33,7'd115}:		p = 14'd3795;
            {7'd33,7'd116}:		p = 14'd3828;
            {7'd33,7'd117}:		p = 14'd3861;
            {7'd33,7'd118}:		p = 14'd3894;
            {7'd33,7'd119}:		p = 14'd3927;
            {7'd33,7'd120}:		p = 14'd3960;
            {7'd33,7'd121}:		p = 14'd3993;
            {7'd33,7'd122}:		p = 14'd4026;
            {7'd33,7'd123}:		p = 14'd4059;
            {7'd33,7'd124}:		p = 14'd4092;
            {7'd33,7'd125}:		p = 14'd4125;
            {7'd33,7'd126}:		p = 14'd4158;
            {7'd33,7'd127}:		p = 14'd4191;
            {7'd34,7'd0}:		p = 14'd0;
            {7'd34,7'd1}:		p = 14'd34;
            {7'd34,7'd2}:		p = 14'd68;
            {7'd34,7'd3}:		p = 14'd102;
            {7'd34,7'd4}:		p = 14'd136;
            {7'd34,7'd5}:		p = 14'd170;
            {7'd34,7'd6}:		p = 14'd204;
            {7'd34,7'd7}:		p = 14'd238;
            {7'd34,7'd8}:		p = 14'd272;
            {7'd34,7'd9}:		p = 14'd306;
            {7'd34,7'd10}:		p = 14'd340;
            {7'd34,7'd11}:		p = 14'd374;
            {7'd34,7'd12}:		p = 14'd408;
            {7'd34,7'd13}:		p = 14'd442;
            {7'd34,7'd14}:		p = 14'd476;
            {7'd34,7'd15}:		p = 14'd510;
            {7'd34,7'd16}:		p = 14'd544;
            {7'd34,7'd17}:		p = 14'd578;
            {7'd34,7'd18}:		p = 14'd612;
            {7'd34,7'd19}:		p = 14'd646;
            {7'd34,7'd20}:		p = 14'd680;
            {7'd34,7'd21}:		p = 14'd714;
            {7'd34,7'd22}:		p = 14'd748;
            {7'd34,7'd23}:		p = 14'd782;
            {7'd34,7'd24}:		p = 14'd816;
            {7'd34,7'd25}:		p = 14'd850;
            {7'd34,7'd26}:		p = 14'd884;
            {7'd34,7'd27}:		p = 14'd918;
            {7'd34,7'd28}:		p = 14'd952;
            {7'd34,7'd29}:		p = 14'd986;
            {7'd34,7'd30}:		p = 14'd1020;
            {7'd34,7'd31}:		p = 14'd1054;
            {7'd34,7'd32}:		p = 14'd1088;
            {7'd34,7'd33}:		p = 14'd1122;
            {7'd34,7'd34}:		p = 14'd1156;
            {7'd34,7'd35}:		p = 14'd1190;
            {7'd34,7'd36}:		p = 14'd1224;
            {7'd34,7'd37}:		p = 14'd1258;
            {7'd34,7'd38}:		p = 14'd1292;
            {7'd34,7'd39}:		p = 14'd1326;
            {7'd34,7'd40}:		p = 14'd1360;
            {7'd34,7'd41}:		p = 14'd1394;
            {7'd34,7'd42}:		p = 14'd1428;
            {7'd34,7'd43}:		p = 14'd1462;
            {7'd34,7'd44}:		p = 14'd1496;
            {7'd34,7'd45}:		p = 14'd1530;
            {7'd34,7'd46}:		p = 14'd1564;
            {7'd34,7'd47}:		p = 14'd1598;
            {7'd34,7'd48}:		p = 14'd1632;
            {7'd34,7'd49}:		p = 14'd1666;
            {7'd34,7'd50}:		p = 14'd1700;
            {7'd34,7'd51}:		p = 14'd1734;
            {7'd34,7'd52}:		p = 14'd1768;
            {7'd34,7'd53}:		p = 14'd1802;
            {7'd34,7'd54}:		p = 14'd1836;
            {7'd34,7'd55}:		p = 14'd1870;
            {7'd34,7'd56}:		p = 14'd1904;
            {7'd34,7'd57}:		p = 14'd1938;
            {7'd34,7'd58}:		p = 14'd1972;
            {7'd34,7'd59}:		p = 14'd2006;
            {7'd34,7'd60}:		p = 14'd2040;
            {7'd34,7'd61}:		p = 14'd2074;
            {7'd34,7'd62}:		p = 14'd2108;
            {7'd34,7'd63}:		p = 14'd2142;
            {7'd34,7'd64}:		p = 14'd2176;
            {7'd34,7'd65}:		p = 14'd2210;
            {7'd34,7'd66}:		p = 14'd2244;
            {7'd34,7'd67}:		p = 14'd2278;
            {7'd34,7'd68}:		p = 14'd2312;
            {7'd34,7'd69}:		p = 14'd2346;
            {7'd34,7'd70}:		p = 14'd2380;
            {7'd34,7'd71}:		p = 14'd2414;
            {7'd34,7'd72}:		p = 14'd2448;
            {7'd34,7'd73}:		p = 14'd2482;
            {7'd34,7'd74}:		p = 14'd2516;
            {7'd34,7'd75}:		p = 14'd2550;
            {7'd34,7'd76}:		p = 14'd2584;
            {7'd34,7'd77}:		p = 14'd2618;
            {7'd34,7'd78}:		p = 14'd2652;
            {7'd34,7'd79}:		p = 14'd2686;
            {7'd34,7'd80}:		p = 14'd2720;
            {7'd34,7'd81}:		p = 14'd2754;
            {7'd34,7'd82}:		p = 14'd2788;
            {7'd34,7'd83}:		p = 14'd2822;
            {7'd34,7'd84}:		p = 14'd2856;
            {7'd34,7'd85}:		p = 14'd2890;
            {7'd34,7'd86}:		p = 14'd2924;
            {7'd34,7'd87}:		p = 14'd2958;
            {7'd34,7'd88}:		p = 14'd2992;
            {7'd34,7'd89}:		p = 14'd3026;
            {7'd34,7'd90}:		p = 14'd3060;
            {7'd34,7'd91}:		p = 14'd3094;
            {7'd34,7'd92}:		p = 14'd3128;
            {7'd34,7'd93}:		p = 14'd3162;
            {7'd34,7'd94}:		p = 14'd3196;
            {7'd34,7'd95}:		p = 14'd3230;
            {7'd34,7'd96}:		p = 14'd3264;
            {7'd34,7'd97}:		p = 14'd3298;
            {7'd34,7'd98}:		p = 14'd3332;
            {7'd34,7'd99}:		p = 14'd3366;
            {7'd34,7'd100}:		p = 14'd3400;
            {7'd34,7'd101}:		p = 14'd3434;
            {7'd34,7'd102}:		p = 14'd3468;
            {7'd34,7'd103}:		p = 14'd3502;
            {7'd34,7'd104}:		p = 14'd3536;
            {7'd34,7'd105}:		p = 14'd3570;
            {7'd34,7'd106}:		p = 14'd3604;
            {7'd34,7'd107}:		p = 14'd3638;
            {7'd34,7'd108}:		p = 14'd3672;
            {7'd34,7'd109}:		p = 14'd3706;
            {7'd34,7'd110}:		p = 14'd3740;
            {7'd34,7'd111}:		p = 14'd3774;
            {7'd34,7'd112}:		p = 14'd3808;
            {7'd34,7'd113}:		p = 14'd3842;
            {7'd34,7'd114}:		p = 14'd3876;
            {7'd34,7'd115}:		p = 14'd3910;
            {7'd34,7'd116}:		p = 14'd3944;
            {7'd34,7'd117}:		p = 14'd3978;
            {7'd34,7'd118}:		p = 14'd4012;
            {7'd34,7'd119}:		p = 14'd4046;
            {7'd34,7'd120}:		p = 14'd4080;
            {7'd34,7'd121}:		p = 14'd4114;
            {7'd34,7'd122}:		p = 14'd4148;
            {7'd34,7'd123}:		p = 14'd4182;
            {7'd34,7'd124}:		p = 14'd4216;
            {7'd34,7'd125}:		p = 14'd4250;
            {7'd34,7'd126}:		p = 14'd4284;
            {7'd34,7'd127}:		p = 14'd4318;
            {7'd35,7'd0}:		p = 14'd0;
            {7'd35,7'd1}:		p = 14'd35;
            {7'd35,7'd2}:		p = 14'd70;
            {7'd35,7'd3}:		p = 14'd105;
            {7'd35,7'd4}:		p = 14'd140;
            {7'd35,7'd5}:		p = 14'd175;
            {7'd35,7'd6}:		p = 14'd210;
            {7'd35,7'd7}:		p = 14'd245;
            {7'd35,7'd8}:		p = 14'd280;
            {7'd35,7'd9}:		p = 14'd315;
            {7'd35,7'd10}:		p = 14'd350;
            {7'd35,7'd11}:		p = 14'd385;
            {7'd35,7'd12}:		p = 14'd420;
            {7'd35,7'd13}:		p = 14'd455;
            {7'd35,7'd14}:		p = 14'd490;
            {7'd35,7'd15}:		p = 14'd525;
            {7'd35,7'd16}:		p = 14'd560;
            {7'd35,7'd17}:		p = 14'd595;
            {7'd35,7'd18}:		p = 14'd630;
            {7'd35,7'd19}:		p = 14'd665;
            {7'd35,7'd20}:		p = 14'd700;
            {7'd35,7'd21}:		p = 14'd735;
            {7'd35,7'd22}:		p = 14'd770;
            {7'd35,7'd23}:		p = 14'd805;
            {7'd35,7'd24}:		p = 14'd840;
            {7'd35,7'd25}:		p = 14'd875;
            {7'd35,7'd26}:		p = 14'd910;
            {7'd35,7'd27}:		p = 14'd945;
            {7'd35,7'd28}:		p = 14'd980;
            {7'd35,7'd29}:		p = 14'd1015;
            {7'd35,7'd30}:		p = 14'd1050;
            {7'd35,7'd31}:		p = 14'd1085;
            {7'd35,7'd32}:		p = 14'd1120;
            {7'd35,7'd33}:		p = 14'd1155;
            {7'd35,7'd34}:		p = 14'd1190;
            {7'd35,7'd35}:		p = 14'd1225;
            {7'd35,7'd36}:		p = 14'd1260;
            {7'd35,7'd37}:		p = 14'd1295;
            {7'd35,7'd38}:		p = 14'd1330;
            {7'd35,7'd39}:		p = 14'd1365;
            {7'd35,7'd40}:		p = 14'd1400;
            {7'd35,7'd41}:		p = 14'd1435;
            {7'd35,7'd42}:		p = 14'd1470;
            {7'd35,7'd43}:		p = 14'd1505;
            {7'd35,7'd44}:		p = 14'd1540;
            {7'd35,7'd45}:		p = 14'd1575;
            {7'd35,7'd46}:		p = 14'd1610;
            {7'd35,7'd47}:		p = 14'd1645;
            {7'd35,7'd48}:		p = 14'd1680;
            {7'd35,7'd49}:		p = 14'd1715;
            {7'd35,7'd50}:		p = 14'd1750;
            {7'd35,7'd51}:		p = 14'd1785;
            {7'd35,7'd52}:		p = 14'd1820;
            {7'd35,7'd53}:		p = 14'd1855;
            {7'd35,7'd54}:		p = 14'd1890;
            {7'd35,7'd55}:		p = 14'd1925;
            {7'd35,7'd56}:		p = 14'd1960;
            {7'd35,7'd57}:		p = 14'd1995;
            {7'd35,7'd58}:		p = 14'd2030;
            {7'd35,7'd59}:		p = 14'd2065;
            {7'd35,7'd60}:		p = 14'd2100;
            {7'd35,7'd61}:		p = 14'd2135;
            {7'd35,7'd62}:		p = 14'd2170;
            {7'd35,7'd63}:		p = 14'd2205;
            {7'd35,7'd64}:		p = 14'd2240;
            {7'd35,7'd65}:		p = 14'd2275;
            {7'd35,7'd66}:		p = 14'd2310;
            {7'd35,7'd67}:		p = 14'd2345;
            {7'd35,7'd68}:		p = 14'd2380;
            {7'd35,7'd69}:		p = 14'd2415;
            {7'd35,7'd70}:		p = 14'd2450;
            {7'd35,7'd71}:		p = 14'd2485;
            {7'd35,7'd72}:		p = 14'd2520;
            {7'd35,7'd73}:		p = 14'd2555;
            {7'd35,7'd74}:		p = 14'd2590;
            {7'd35,7'd75}:		p = 14'd2625;
            {7'd35,7'd76}:		p = 14'd2660;
            {7'd35,7'd77}:		p = 14'd2695;
            {7'd35,7'd78}:		p = 14'd2730;
            {7'd35,7'd79}:		p = 14'd2765;
            {7'd35,7'd80}:		p = 14'd2800;
            {7'd35,7'd81}:		p = 14'd2835;
            {7'd35,7'd82}:		p = 14'd2870;
            {7'd35,7'd83}:		p = 14'd2905;
            {7'd35,7'd84}:		p = 14'd2940;
            {7'd35,7'd85}:		p = 14'd2975;
            {7'd35,7'd86}:		p = 14'd3010;
            {7'd35,7'd87}:		p = 14'd3045;
            {7'd35,7'd88}:		p = 14'd3080;
            {7'd35,7'd89}:		p = 14'd3115;
            {7'd35,7'd90}:		p = 14'd3150;
            {7'd35,7'd91}:		p = 14'd3185;
            {7'd35,7'd92}:		p = 14'd3220;
            {7'd35,7'd93}:		p = 14'd3255;
            {7'd35,7'd94}:		p = 14'd3290;
            {7'd35,7'd95}:		p = 14'd3325;
            {7'd35,7'd96}:		p = 14'd3360;
            {7'd35,7'd97}:		p = 14'd3395;
            {7'd35,7'd98}:		p = 14'd3430;
            {7'd35,7'd99}:		p = 14'd3465;
            {7'd35,7'd100}:		p = 14'd3500;
            {7'd35,7'd101}:		p = 14'd3535;
            {7'd35,7'd102}:		p = 14'd3570;
            {7'd35,7'd103}:		p = 14'd3605;
            {7'd35,7'd104}:		p = 14'd3640;
            {7'd35,7'd105}:		p = 14'd3675;
            {7'd35,7'd106}:		p = 14'd3710;
            {7'd35,7'd107}:		p = 14'd3745;
            {7'd35,7'd108}:		p = 14'd3780;
            {7'd35,7'd109}:		p = 14'd3815;
            {7'd35,7'd110}:		p = 14'd3850;
            {7'd35,7'd111}:		p = 14'd3885;
            {7'd35,7'd112}:		p = 14'd3920;
            {7'd35,7'd113}:		p = 14'd3955;
            {7'd35,7'd114}:		p = 14'd3990;
            {7'd35,7'd115}:		p = 14'd4025;
            {7'd35,7'd116}:		p = 14'd4060;
            {7'd35,7'd117}:		p = 14'd4095;
            {7'd35,7'd118}:		p = 14'd4130;
            {7'd35,7'd119}:		p = 14'd4165;
            {7'd35,7'd120}:		p = 14'd4200;
            {7'd35,7'd121}:		p = 14'd4235;
            {7'd35,7'd122}:		p = 14'd4270;
            {7'd35,7'd123}:		p = 14'd4305;
            {7'd35,7'd124}:		p = 14'd4340;
            {7'd35,7'd125}:		p = 14'd4375;
            {7'd35,7'd126}:		p = 14'd4410;
            {7'd35,7'd127}:		p = 14'd4445;
            {7'd36,7'd0}:		p = 14'd0;
            {7'd36,7'd1}:		p = 14'd36;
            {7'd36,7'd2}:		p = 14'd72;
            {7'd36,7'd3}:		p = 14'd108;
            {7'd36,7'd4}:		p = 14'd144;
            {7'd36,7'd5}:		p = 14'd180;
            {7'd36,7'd6}:		p = 14'd216;
            {7'd36,7'd7}:		p = 14'd252;
            {7'd36,7'd8}:		p = 14'd288;
            {7'd36,7'd9}:		p = 14'd324;
            {7'd36,7'd10}:		p = 14'd360;
            {7'd36,7'd11}:		p = 14'd396;
            {7'd36,7'd12}:		p = 14'd432;
            {7'd36,7'd13}:		p = 14'd468;
            {7'd36,7'd14}:		p = 14'd504;
            {7'd36,7'd15}:		p = 14'd540;
            {7'd36,7'd16}:		p = 14'd576;
            {7'd36,7'd17}:		p = 14'd612;
            {7'd36,7'd18}:		p = 14'd648;
            {7'd36,7'd19}:		p = 14'd684;
            {7'd36,7'd20}:		p = 14'd720;
            {7'd36,7'd21}:		p = 14'd756;
            {7'd36,7'd22}:		p = 14'd792;
            {7'd36,7'd23}:		p = 14'd828;
            {7'd36,7'd24}:		p = 14'd864;
            {7'd36,7'd25}:		p = 14'd900;
            {7'd36,7'd26}:		p = 14'd936;
            {7'd36,7'd27}:		p = 14'd972;
            {7'd36,7'd28}:		p = 14'd1008;
            {7'd36,7'd29}:		p = 14'd1044;
            {7'd36,7'd30}:		p = 14'd1080;
            {7'd36,7'd31}:		p = 14'd1116;
            {7'd36,7'd32}:		p = 14'd1152;
            {7'd36,7'd33}:		p = 14'd1188;
            {7'd36,7'd34}:		p = 14'd1224;
            {7'd36,7'd35}:		p = 14'd1260;
            {7'd36,7'd36}:		p = 14'd1296;
            {7'd36,7'd37}:		p = 14'd1332;
            {7'd36,7'd38}:		p = 14'd1368;
            {7'd36,7'd39}:		p = 14'd1404;
            {7'd36,7'd40}:		p = 14'd1440;
            {7'd36,7'd41}:		p = 14'd1476;
            {7'd36,7'd42}:		p = 14'd1512;
            {7'd36,7'd43}:		p = 14'd1548;
            {7'd36,7'd44}:		p = 14'd1584;
            {7'd36,7'd45}:		p = 14'd1620;
            {7'd36,7'd46}:		p = 14'd1656;
            {7'd36,7'd47}:		p = 14'd1692;
            {7'd36,7'd48}:		p = 14'd1728;
            {7'd36,7'd49}:		p = 14'd1764;
            {7'd36,7'd50}:		p = 14'd1800;
            {7'd36,7'd51}:		p = 14'd1836;
            {7'd36,7'd52}:		p = 14'd1872;
            {7'd36,7'd53}:		p = 14'd1908;
            {7'd36,7'd54}:		p = 14'd1944;
            {7'd36,7'd55}:		p = 14'd1980;
            {7'd36,7'd56}:		p = 14'd2016;
            {7'd36,7'd57}:		p = 14'd2052;
            {7'd36,7'd58}:		p = 14'd2088;
            {7'd36,7'd59}:		p = 14'd2124;
            {7'd36,7'd60}:		p = 14'd2160;
            {7'd36,7'd61}:		p = 14'd2196;
            {7'd36,7'd62}:		p = 14'd2232;
            {7'd36,7'd63}:		p = 14'd2268;
            {7'd36,7'd64}:		p = 14'd2304;
            {7'd36,7'd65}:		p = 14'd2340;
            {7'd36,7'd66}:		p = 14'd2376;
            {7'd36,7'd67}:		p = 14'd2412;
            {7'd36,7'd68}:		p = 14'd2448;
            {7'd36,7'd69}:		p = 14'd2484;
            {7'd36,7'd70}:		p = 14'd2520;
            {7'd36,7'd71}:		p = 14'd2556;
            {7'd36,7'd72}:		p = 14'd2592;
            {7'd36,7'd73}:		p = 14'd2628;
            {7'd36,7'd74}:		p = 14'd2664;
            {7'd36,7'd75}:		p = 14'd2700;
            {7'd36,7'd76}:		p = 14'd2736;
            {7'd36,7'd77}:		p = 14'd2772;
            {7'd36,7'd78}:		p = 14'd2808;
            {7'd36,7'd79}:		p = 14'd2844;
            {7'd36,7'd80}:		p = 14'd2880;
            {7'd36,7'd81}:		p = 14'd2916;
            {7'd36,7'd82}:		p = 14'd2952;
            {7'd36,7'd83}:		p = 14'd2988;
            {7'd36,7'd84}:		p = 14'd3024;
            {7'd36,7'd85}:		p = 14'd3060;
            {7'd36,7'd86}:		p = 14'd3096;
            {7'd36,7'd87}:		p = 14'd3132;
            {7'd36,7'd88}:		p = 14'd3168;
            {7'd36,7'd89}:		p = 14'd3204;
            {7'd36,7'd90}:		p = 14'd3240;
            {7'd36,7'd91}:		p = 14'd3276;
            {7'd36,7'd92}:		p = 14'd3312;
            {7'd36,7'd93}:		p = 14'd3348;
            {7'd36,7'd94}:		p = 14'd3384;
            {7'd36,7'd95}:		p = 14'd3420;
            {7'd36,7'd96}:		p = 14'd3456;
            {7'd36,7'd97}:		p = 14'd3492;
            {7'd36,7'd98}:		p = 14'd3528;
            {7'd36,7'd99}:		p = 14'd3564;
            {7'd36,7'd100}:		p = 14'd3600;
            {7'd36,7'd101}:		p = 14'd3636;
            {7'd36,7'd102}:		p = 14'd3672;
            {7'd36,7'd103}:		p = 14'd3708;
            {7'd36,7'd104}:		p = 14'd3744;
            {7'd36,7'd105}:		p = 14'd3780;
            {7'd36,7'd106}:		p = 14'd3816;
            {7'd36,7'd107}:		p = 14'd3852;
            {7'd36,7'd108}:		p = 14'd3888;
            {7'd36,7'd109}:		p = 14'd3924;
            {7'd36,7'd110}:		p = 14'd3960;
            {7'd36,7'd111}:		p = 14'd3996;
            {7'd36,7'd112}:		p = 14'd4032;
            {7'd36,7'd113}:		p = 14'd4068;
            {7'd36,7'd114}:		p = 14'd4104;
            {7'd36,7'd115}:		p = 14'd4140;
            {7'd36,7'd116}:		p = 14'd4176;
            {7'd36,7'd117}:		p = 14'd4212;
            {7'd36,7'd118}:		p = 14'd4248;
            {7'd36,7'd119}:		p = 14'd4284;
            {7'd36,7'd120}:		p = 14'd4320;
            {7'd36,7'd121}:		p = 14'd4356;
            {7'd36,7'd122}:		p = 14'd4392;
            {7'd36,7'd123}:		p = 14'd4428;
            {7'd36,7'd124}:		p = 14'd4464;
            {7'd36,7'd125}:		p = 14'd4500;
            {7'd36,7'd126}:		p = 14'd4536;
            {7'd36,7'd127}:		p = 14'd4572;
            {7'd37,7'd0}:		p = 14'd0;
            {7'd37,7'd1}:		p = 14'd37;
            {7'd37,7'd2}:		p = 14'd74;
            {7'd37,7'd3}:		p = 14'd111;
            {7'd37,7'd4}:		p = 14'd148;
            {7'd37,7'd5}:		p = 14'd185;
            {7'd37,7'd6}:		p = 14'd222;
            {7'd37,7'd7}:		p = 14'd259;
            {7'd37,7'd8}:		p = 14'd296;
            {7'd37,7'd9}:		p = 14'd333;
            {7'd37,7'd10}:		p = 14'd370;
            {7'd37,7'd11}:		p = 14'd407;
            {7'd37,7'd12}:		p = 14'd444;
            {7'd37,7'd13}:		p = 14'd481;
            {7'd37,7'd14}:		p = 14'd518;
            {7'd37,7'd15}:		p = 14'd555;
            {7'd37,7'd16}:		p = 14'd592;
            {7'd37,7'd17}:		p = 14'd629;
            {7'd37,7'd18}:		p = 14'd666;
            {7'd37,7'd19}:		p = 14'd703;
            {7'd37,7'd20}:		p = 14'd740;
            {7'd37,7'd21}:		p = 14'd777;
            {7'd37,7'd22}:		p = 14'd814;
            {7'd37,7'd23}:		p = 14'd851;
            {7'd37,7'd24}:		p = 14'd888;
            {7'd37,7'd25}:		p = 14'd925;
            {7'd37,7'd26}:		p = 14'd962;
            {7'd37,7'd27}:		p = 14'd999;
            {7'd37,7'd28}:		p = 14'd1036;
            {7'd37,7'd29}:		p = 14'd1073;
            {7'd37,7'd30}:		p = 14'd1110;
            {7'd37,7'd31}:		p = 14'd1147;
            {7'd37,7'd32}:		p = 14'd1184;
            {7'd37,7'd33}:		p = 14'd1221;
            {7'd37,7'd34}:		p = 14'd1258;
            {7'd37,7'd35}:		p = 14'd1295;
            {7'd37,7'd36}:		p = 14'd1332;
            {7'd37,7'd37}:		p = 14'd1369;
            {7'd37,7'd38}:		p = 14'd1406;
            {7'd37,7'd39}:		p = 14'd1443;
            {7'd37,7'd40}:		p = 14'd1480;
            {7'd37,7'd41}:		p = 14'd1517;
            {7'd37,7'd42}:		p = 14'd1554;
            {7'd37,7'd43}:		p = 14'd1591;
            {7'd37,7'd44}:		p = 14'd1628;
            {7'd37,7'd45}:		p = 14'd1665;
            {7'd37,7'd46}:		p = 14'd1702;
            {7'd37,7'd47}:		p = 14'd1739;
            {7'd37,7'd48}:		p = 14'd1776;
            {7'd37,7'd49}:		p = 14'd1813;
            {7'd37,7'd50}:		p = 14'd1850;
            {7'd37,7'd51}:		p = 14'd1887;
            {7'd37,7'd52}:		p = 14'd1924;
            {7'd37,7'd53}:		p = 14'd1961;
            {7'd37,7'd54}:		p = 14'd1998;
            {7'd37,7'd55}:		p = 14'd2035;
            {7'd37,7'd56}:		p = 14'd2072;
            {7'd37,7'd57}:		p = 14'd2109;
            {7'd37,7'd58}:		p = 14'd2146;
            {7'd37,7'd59}:		p = 14'd2183;
            {7'd37,7'd60}:		p = 14'd2220;
            {7'd37,7'd61}:		p = 14'd2257;
            {7'd37,7'd62}:		p = 14'd2294;
            {7'd37,7'd63}:		p = 14'd2331;
            {7'd37,7'd64}:		p = 14'd2368;
            {7'd37,7'd65}:		p = 14'd2405;
            {7'd37,7'd66}:		p = 14'd2442;
            {7'd37,7'd67}:		p = 14'd2479;
            {7'd37,7'd68}:		p = 14'd2516;
            {7'd37,7'd69}:		p = 14'd2553;
            {7'd37,7'd70}:		p = 14'd2590;
            {7'd37,7'd71}:		p = 14'd2627;
            {7'd37,7'd72}:		p = 14'd2664;
            {7'd37,7'd73}:		p = 14'd2701;
            {7'd37,7'd74}:		p = 14'd2738;
            {7'd37,7'd75}:		p = 14'd2775;
            {7'd37,7'd76}:		p = 14'd2812;
            {7'd37,7'd77}:		p = 14'd2849;
            {7'd37,7'd78}:		p = 14'd2886;
            {7'd37,7'd79}:		p = 14'd2923;
            {7'd37,7'd80}:		p = 14'd2960;
            {7'd37,7'd81}:		p = 14'd2997;
            {7'd37,7'd82}:		p = 14'd3034;
            {7'd37,7'd83}:		p = 14'd3071;
            {7'd37,7'd84}:		p = 14'd3108;
            {7'd37,7'd85}:		p = 14'd3145;
            {7'd37,7'd86}:		p = 14'd3182;
            {7'd37,7'd87}:		p = 14'd3219;
            {7'd37,7'd88}:		p = 14'd3256;
            {7'd37,7'd89}:		p = 14'd3293;
            {7'd37,7'd90}:		p = 14'd3330;
            {7'd37,7'd91}:		p = 14'd3367;
            {7'd37,7'd92}:		p = 14'd3404;
            {7'd37,7'd93}:		p = 14'd3441;
            {7'd37,7'd94}:		p = 14'd3478;
            {7'd37,7'd95}:		p = 14'd3515;
            {7'd37,7'd96}:		p = 14'd3552;
            {7'd37,7'd97}:		p = 14'd3589;
            {7'd37,7'd98}:		p = 14'd3626;
            {7'd37,7'd99}:		p = 14'd3663;
            {7'd37,7'd100}:		p = 14'd3700;
            {7'd37,7'd101}:		p = 14'd3737;
            {7'd37,7'd102}:		p = 14'd3774;
            {7'd37,7'd103}:		p = 14'd3811;
            {7'd37,7'd104}:		p = 14'd3848;
            {7'd37,7'd105}:		p = 14'd3885;
            {7'd37,7'd106}:		p = 14'd3922;
            {7'd37,7'd107}:		p = 14'd3959;
            {7'd37,7'd108}:		p = 14'd3996;
            {7'd37,7'd109}:		p = 14'd4033;
            {7'd37,7'd110}:		p = 14'd4070;
            {7'd37,7'd111}:		p = 14'd4107;
            {7'd37,7'd112}:		p = 14'd4144;
            {7'd37,7'd113}:		p = 14'd4181;
            {7'd37,7'd114}:		p = 14'd4218;
            {7'd37,7'd115}:		p = 14'd4255;
            {7'd37,7'd116}:		p = 14'd4292;
            {7'd37,7'd117}:		p = 14'd4329;
            {7'd37,7'd118}:		p = 14'd4366;
            {7'd37,7'd119}:		p = 14'd4403;
            {7'd37,7'd120}:		p = 14'd4440;
            {7'd37,7'd121}:		p = 14'd4477;
            {7'd37,7'd122}:		p = 14'd4514;
            {7'd37,7'd123}:		p = 14'd4551;
            {7'd37,7'd124}:		p = 14'd4588;
            {7'd37,7'd125}:		p = 14'd4625;
            {7'd37,7'd126}:		p = 14'd4662;
            {7'd37,7'd127}:		p = 14'd4699;
            {7'd38,7'd0}:		p = 14'd0;
            {7'd38,7'd1}:		p = 14'd38;
            {7'd38,7'd2}:		p = 14'd76;
            {7'd38,7'd3}:		p = 14'd114;
            {7'd38,7'd4}:		p = 14'd152;
            {7'd38,7'd5}:		p = 14'd190;
            {7'd38,7'd6}:		p = 14'd228;
            {7'd38,7'd7}:		p = 14'd266;
            {7'd38,7'd8}:		p = 14'd304;
            {7'd38,7'd9}:		p = 14'd342;
            {7'd38,7'd10}:		p = 14'd380;
            {7'd38,7'd11}:		p = 14'd418;
            {7'd38,7'd12}:		p = 14'd456;
            {7'd38,7'd13}:		p = 14'd494;
            {7'd38,7'd14}:		p = 14'd532;
            {7'd38,7'd15}:		p = 14'd570;
            {7'd38,7'd16}:		p = 14'd608;
            {7'd38,7'd17}:		p = 14'd646;
            {7'd38,7'd18}:		p = 14'd684;
            {7'd38,7'd19}:		p = 14'd722;
            {7'd38,7'd20}:		p = 14'd760;
            {7'd38,7'd21}:		p = 14'd798;
            {7'd38,7'd22}:		p = 14'd836;
            {7'd38,7'd23}:		p = 14'd874;
            {7'd38,7'd24}:		p = 14'd912;
            {7'd38,7'd25}:		p = 14'd950;
            {7'd38,7'd26}:		p = 14'd988;
            {7'd38,7'd27}:		p = 14'd1026;
            {7'd38,7'd28}:		p = 14'd1064;
            {7'd38,7'd29}:		p = 14'd1102;
            {7'd38,7'd30}:		p = 14'd1140;
            {7'd38,7'd31}:		p = 14'd1178;
            {7'd38,7'd32}:		p = 14'd1216;
            {7'd38,7'd33}:		p = 14'd1254;
            {7'd38,7'd34}:		p = 14'd1292;
            {7'd38,7'd35}:		p = 14'd1330;
            {7'd38,7'd36}:		p = 14'd1368;
            {7'd38,7'd37}:		p = 14'd1406;
            {7'd38,7'd38}:		p = 14'd1444;
            {7'd38,7'd39}:		p = 14'd1482;
            {7'd38,7'd40}:		p = 14'd1520;
            {7'd38,7'd41}:		p = 14'd1558;
            {7'd38,7'd42}:		p = 14'd1596;
            {7'd38,7'd43}:		p = 14'd1634;
            {7'd38,7'd44}:		p = 14'd1672;
            {7'd38,7'd45}:		p = 14'd1710;
            {7'd38,7'd46}:		p = 14'd1748;
            {7'd38,7'd47}:		p = 14'd1786;
            {7'd38,7'd48}:		p = 14'd1824;
            {7'd38,7'd49}:		p = 14'd1862;
            {7'd38,7'd50}:		p = 14'd1900;
            {7'd38,7'd51}:		p = 14'd1938;
            {7'd38,7'd52}:		p = 14'd1976;
            {7'd38,7'd53}:		p = 14'd2014;
            {7'd38,7'd54}:		p = 14'd2052;
            {7'd38,7'd55}:		p = 14'd2090;
            {7'd38,7'd56}:		p = 14'd2128;
            {7'd38,7'd57}:		p = 14'd2166;
            {7'd38,7'd58}:		p = 14'd2204;
            {7'd38,7'd59}:		p = 14'd2242;
            {7'd38,7'd60}:		p = 14'd2280;
            {7'd38,7'd61}:		p = 14'd2318;
            {7'd38,7'd62}:		p = 14'd2356;
            {7'd38,7'd63}:		p = 14'd2394;
            {7'd38,7'd64}:		p = 14'd2432;
            {7'd38,7'd65}:		p = 14'd2470;
            {7'd38,7'd66}:		p = 14'd2508;
            {7'd38,7'd67}:		p = 14'd2546;
            {7'd38,7'd68}:		p = 14'd2584;
            {7'd38,7'd69}:		p = 14'd2622;
            {7'd38,7'd70}:		p = 14'd2660;
            {7'd38,7'd71}:		p = 14'd2698;
            {7'd38,7'd72}:		p = 14'd2736;
            {7'd38,7'd73}:		p = 14'd2774;
            {7'd38,7'd74}:		p = 14'd2812;
            {7'd38,7'd75}:		p = 14'd2850;
            {7'd38,7'd76}:		p = 14'd2888;
            {7'd38,7'd77}:		p = 14'd2926;
            {7'd38,7'd78}:		p = 14'd2964;
            {7'd38,7'd79}:		p = 14'd3002;
            {7'd38,7'd80}:		p = 14'd3040;
            {7'd38,7'd81}:		p = 14'd3078;
            {7'd38,7'd82}:		p = 14'd3116;
            {7'd38,7'd83}:		p = 14'd3154;
            {7'd38,7'd84}:		p = 14'd3192;
            {7'd38,7'd85}:		p = 14'd3230;
            {7'd38,7'd86}:		p = 14'd3268;
            {7'd38,7'd87}:		p = 14'd3306;
            {7'd38,7'd88}:		p = 14'd3344;
            {7'd38,7'd89}:		p = 14'd3382;
            {7'd38,7'd90}:		p = 14'd3420;
            {7'd38,7'd91}:		p = 14'd3458;
            {7'd38,7'd92}:		p = 14'd3496;
            {7'd38,7'd93}:		p = 14'd3534;
            {7'd38,7'd94}:		p = 14'd3572;
            {7'd38,7'd95}:		p = 14'd3610;
            {7'd38,7'd96}:		p = 14'd3648;
            {7'd38,7'd97}:		p = 14'd3686;
            {7'd38,7'd98}:		p = 14'd3724;
            {7'd38,7'd99}:		p = 14'd3762;
            {7'd38,7'd100}:		p = 14'd3800;
            {7'd38,7'd101}:		p = 14'd3838;
            {7'd38,7'd102}:		p = 14'd3876;
            {7'd38,7'd103}:		p = 14'd3914;
            {7'd38,7'd104}:		p = 14'd3952;
            {7'd38,7'd105}:		p = 14'd3990;
            {7'd38,7'd106}:		p = 14'd4028;
            {7'd38,7'd107}:		p = 14'd4066;
            {7'd38,7'd108}:		p = 14'd4104;
            {7'd38,7'd109}:		p = 14'd4142;
            {7'd38,7'd110}:		p = 14'd4180;
            {7'd38,7'd111}:		p = 14'd4218;
            {7'd38,7'd112}:		p = 14'd4256;
            {7'd38,7'd113}:		p = 14'd4294;
            {7'd38,7'd114}:		p = 14'd4332;
            {7'd38,7'd115}:		p = 14'd4370;
            {7'd38,7'd116}:		p = 14'd4408;
            {7'd38,7'd117}:		p = 14'd4446;
            {7'd38,7'd118}:		p = 14'd4484;
            {7'd38,7'd119}:		p = 14'd4522;
            {7'd38,7'd120}:		p = 14'd4560;
            {7'd38,7'd121}:		p = 14'd4598;
            {7'd38,7'd122}:		p = 14'd4636;
            {7'd38,7'd123}:		p = 14'd4674;
            {7'd38,7'd124}:		p = 14'd4712;
            {7'd38,7'd125}:		p = 14'd4750;
            {7'd38,7'd126}:		p = 14'd4788;
            {7'd38,7'd127}:		p = 14'd4826;
            {7'd39,7'd0}:		p = 14'd0;
            {7'd39,7'd1}:		p = 14'd39;
            {7'd39,7'd2}:		p = 14'd78;
            {7'd39,7'd3}:		p = 14'd117;
            {7'd39,7'd4}:		p = 14'd156;
            {7'd39,7'd5}:		p = 14'd195;
            {7'd39,7'd6}:		p = 14'd234;
            {7'd39,7'd7}:		p = 14'd273;
            {7'd39,7'd8}:		p = 14'd312;
            {7'd39,7'd9}:		p = 14'd351;
            {7'd39,7'd10}:		p = 14'd390;
            {7'd39,7'd11}:		p = 14'd429;
            {7'd39,7'd12}:		p = 14'd468;
            {7'd39,7'd13}:		p = 14'd507;
            {7'd39,7'd14}:		p = 14'd546;
            {7'd39,7'd15}:		p = 14'd585;
            {7'd39,7'd16}:		p = 14'd624;
            {7'd39,7'd17}:		p = 14'd663;
            {7'd39,7'd18}:		p = 14'd702;
            {7'd39,7'd19}:		p = 14'd741;
            {7'd39,7'd20}:		p = 14'd780;
            {7'd39,7'd21}:		p = 14'd819;
            {7'd39,7'd22}:		p = 14'd858;
            {7'd39,7'd23}:		p = 14'd897;
            {7'd39,7'd24}:		p = 14'd936;
            {7'd39,7'd25}:		p = 14'd975;
            {7'd39,7'd26}:		p = 14'd1014;
            {7'd39,7'd27}:		p = 14'd1053;
            {7'd39,7'd28}:		p = 14'd1092;
            {7'd39,7'd29}:		p = 14'd1131;
            {7'd39,7'd30}:		p = 14'd1170;
            {7'd39,7'd31}:		p = 14'd1209;
            {7'd39,7'd32}:		p = 14'd1248;
            {7'd39,7'd33}:		p = 14'd1287;
            {7'd39,7'd34}:		p = 14'd1326;
            {7'd39,7'd35}:		p = 14'd1365;
            {7'd39,7'd36}:		p = 14'd1404;
            {7'd39,7'd37}:		p = 14'd1443;
            {7'd39,7'd38}:		p = 14'd1482;
            {7'd39,7'd39}:		p = 14'd1521;
            {7'd39,7'd40}:		p = 14'd1560;
            {7'd39,7'd41}:		p = 14'd1599;
            {7'd39,7'd42}:		p = 14'd1638;
            {7'd39,7'd43}:		p = 14'd1677;
            {7'd39,7'd44}:		p = 14'd1716;
            {7'd39,7'd45}:		p = 14'd1755;
            {7'd39,7'd46}:		p = 14'd1794;
            {7'd39,7'd47}:		p = 14'd1833;
            {7'd39,7'd48}:		p = 14'd1872;
            {7'd39,7'd49}:		p = 14'd1911;
            {7'd39,7'd50}:		p = 14'd1950;
            {7'd39,7'd51}:		p = 14'd1989;
            {7'd39,7'd52}:		p = 14'd2028;
            {7'd39,7'd53}:		p = 14'd2067;
            {7'd39,7'd54}:		p = 14'd2106;
            {7'd39,7'd55}:		p = 14'd2145;
            {7'd39,7'd56}:		p = 14'd2184;
            {7'd39,7'd57}:		p = 14'd2223;
            {7'd39,7'd58}:		p = 14'd2262;
            {7'd39,7'd59}:		p = 14'd2301;
            {7'd39,7'd60}:		p = 14'd2340;
            {7'd39,7'd61}:		p = 14'd2379;
            {7'd39,7'd62}:		p = 14'd2418;
            {7'd39,7'd63}:		p = 14'd2457;
            {7'd39,7'd64}:		p = 14'd2496;
            {7'd39,7'd65}:		p = 14'd2535;
            {7'd39,7'd66}:		p = 14'd2574;
            {7'd39,7'd67}:		p = 14'd2613;
            {7'd39,7'd68}:		p = 14'd2652;
            {7'd39,7'd69}:		p = 14'd2691;
            {7'd39,7'd70}:		p = 14'd2730;
            {7'd39,7'd71}:		p = 14'd2769;
            {7'd39,7'd72}:		p = 14'd2808;
            {7'd39,7'd73}:		p = 14'd2847;
            {7'd39,7'd74}:		p = 14'd2886;
            {7'd39,7'd75}:		p = 14'd2925;
            {7'd39,7'd76}:		p = 14'd2964;
            {7'd39,7'd77}:		p = 14'd3003;
            {7'd39,7'd78}:		p = 14'd3042;
            {7'd39,7'd79}:		p = 14'd3081;
            {7'd39,7'd80}:		p = 14'd3120;
            {7'd39,7'd81}:		p = 14'd3159;
            {7'd39,7'd82}:		p = 14'd3198;
            {7'd39,7'd83}:		p = 14'd3237;
            {7'd39,7'd84}:		p = 14'd3276;
            {7'd39,7'd85}:		p = 14'd3315;
            {7'd39,7'd86}:		p = 14'd3354;
            {7'd39,7'd87}:		p = 14'd3393;
            {7'd39,7'd88}:		p = 14'd3432;
            {7'd39,7'd89}:		p = 14'd3471;
            {7'd39,7'd90}:		p = 14'd3510;
            {7'd39,7'd91}:		p = 14'd3549;
            {7'd39,7'd92}:		p = 14'd3588;
            {7'd39,7'd93}:		p = 14'd3627;
            {7'd39,7'd94}:		p = 14'd3666;
            {7'd39,7'd95}:		p = 14'd3705;
            {7'd39,7'd96}:		p = 14'd3744;
            {7'd39,7'd97}:		p = 14'd3783;
            {7'd39,7'd98}:		p = 14'd3822;
            {7'd39,7'd99}:		p = 14'd3861;
            {7'd39,7'd100}:		p = 14'd3900;
            {7'd39,7'd101}:		p = 14'd3939;
            {7'd39,7'd102}:		p = 14'd3978;
            {7'd39,7'd103}:		p = 14'd4017;
            {7'd39,7'd104}:		p = 14'd4056;
            {7'd39,7'd105}:		p = 14'd4095;
            {7'd39,7'd106}:		p = 14'd4134;
            {7'd39,7'd107}:		p = 14'd4173;
            {7'd39,7'd108}:		p = 14'd4212;
            {7'd39,7'd109}:		p = 14'd4251;
            {7'd39,7'd110}:		p = 14'd4290;
            {7'd39,7'd111}:		p = 14'd4329;
            {7'd39,7'd112}:		p = 14'd4368;
            {7'd39,7'd113}:		p = 14'd4407;
            {7'd39,7'd114}:		p = 14'd4446;
            {7'd39,7'd115}:		p = 14'd4485;
            {7'd39,7'd116}:		p = 14'd4524;
            {7'd39,7'd117}:		p = 14'd4563;
            {7'd39,7'd118}:		p = 14'd4602;
            {7'd39,7'd119}:		p = 14'd4641;
            {7'd39,7'd120}:		p = 14'd4680;
            {7'd39,7'd121}:		p = 14'd4719;
            {7'd39,7'd122}:		p = 14'd4758;
            {7'd39,7'd123}:		p = 14'd4797;
            {7'd39,7'd124}:		p = 14'd4836;
            {7'd39,7'd125}:		p = 14'd4875;
            {7'd39,7'd126}:		p = 14'd4914;
            {7'd39,7'd127}:		p = 14'd4953;
            {7'd40,7'd0}:		p = 14'd0;
            {7'd40,7'd1}:		p = 14'd40;
            {7'd40,7'd2}:		p = 14'd80;
            {7'd40,7'd3}:		p = 14'd120;
            {7'd40,7'd4}:		p = 14'd160;
            {7'd40,7'd5}:		p = 14'd200;
            {7'd40,7'd6}:		p = 14'd240;
            {7'd40,7'd7}:		p = 14'd280;
            {7'd40,7'd8}:		p = 14'd320;
            {7'd40,7'd9}:		p = 14'd360;
            {7'd40,7'd10}:		p = 14'd400;
            {7'd40,7'd11}:		p = 14'd440;
            {7'd40,7'd12}:		p = 14'd480;
            {7'd40,7'd13}:		p = 14'd520;
            {7'd40,7'd14}:		p = 14'd560;
            {7'd40,7'd15}:		p = 14'd600;
            {7'd40,7'd16}:		p = 14'd640;
            {7'd40,7'd17}:		p = 14'd680;
            {7'd40,7'd18}:		p = 14'd720;
            {7'd40,7'd19}:		p = 14'd760;
            {7'd40,7'd20}:		p = 14'd800;
            {7'd40,7'd21}:		p = 14'd840;
            {7'd40,7'd22}:		p = 14'd880;
            {7'd40,7'd23}:		p = 14'd920;
            {7'd40,7'd24}:		p = 14'd960;
            {7'd40,7'd25}:		p = 14'd1000;
            {7'd40,7'd26}:		p = 14'd1040;
            {7'd40,7'd27}:		p = 14'd1080;
            {7'd40,7'd28}:		p = 14'd1120;
            {7'd40,7'd29}:		p = 14'd1160;
            {7'd40,7'd30}:		p = 14'd1200;
            {7'd40,7'd31}:		p = 14'd1240;
            {7'd40,7'd32}:		p = 14'd1280;
            {7'd40,7'd33}:		p = 14'd1320;
            {7'd40,7'd34}:		p = 14'd1360;
            {7'd40,7'd35}:		p = 14'd1400;
            {7'd40,7'd36}:		p = 14'd1440;
            {7'd40,7'd37}:		p = 14'd1480;
            {7'd40,7'd38}:		p = 14'd1520;
            {7'd40,7'd39}:		p = 14'd1560;
            {7'd40,7'd40}:		p = 14'd1600;
            {7'd40,7'd41}:		p = 14'd1640;
            {7'd40,7'd42}:		p = 14'd1680;
            {7'd40,7'd43}:		p = 14'd1720;
            {7'd40,7'd44}:		p = 14'd1760;
            {7'd40,7'd45}:		p = 14'd1800;
            {7'd40,7'd46}:		p = 14'd1840;
            {7'd40,7'd47}:		p = 14'd1880;
            {7'd40,7'd48}:		p = 14'd1920;
            {7'd40,7'd49}:		p = 14'd1960;
            {7'd40,7'd50}:		p = 14'd2000;
            {7'd40,7'd51}:		p = 14'd2040;
            {7'd40,7'd52}:		p = 14'd2080;
            {7'd40,7'd53}:		p = 14'd2120;
            {7'd40,7'd54}:		p = 14'd2160;
            {7'd40,7'd55}:		p = 14'd2200;
            {7'd40,7'd56}:		p = 14'd2240;
            {7'd40,7'd57}:		p = 14'd2280;
            {7'd40,7'd58}:		p = 14'd2320;
            {7'd40,7'd59}:		p = 14'd2360;
            {7'd40,7'd60}:		p = 14'd2400;
            {7'd40,7'd61}:		p = 14'd2440;
            {7'd40,7'd62}:		p = 14'd2480;
            {7'd40,7'd63}:		p = 14'd2520;
            {7'd40,7'd64}:		p = 14'd2560;
            {7'd40,7'd65}:		p = 14'd2600;
            {7'd40,7'd66}:		p = 14'd2640;
            {7'd40,7'd67}:		p = 14'd2680;
            {7'd40,7'd68}:		p = 14'd2720;
            {7'd40,7'd69}:		p = 14'd2760;
            {7'd40,7'd70}:		p = 14'd2800;
            {7'd40,7'd71}:		p = 14'd2840;
            {7'd40,7'd72}:		p = 14'd2880;
            {7'd40,7'd73}:		p = 14'd2920;
            {7'd40,7'd74}:		p = 14'd2960;
            {7'd40,7'd75}:		p = 14'd3000;
            {7'd40,7'd76}:		p = 14'd3040;
            {7'd40,7'd77}:		p = 14'd3080;
            {7'd40,7'd78}:		p = 14'd3120;
            {7'd40,7'd79}:		p = 14'd3160;
            {7'd40,7'd80}:		p = 14'd3200;
            {7'd40,7'd81}:		p = 14'd3240;
            {7'd40,7'd82}:		p = 14'd3280;
            {7'd40,7'd83}:		p = 14'd3320;
            {7'd40,7'd84}:		p = 14'd3360;
            {7'd40,7'd85}:		p = 14'd3400;
            {7'd40,7'd86}:		p = 14'd3440;
            {7'd40,7'd87}:		p = 14'd3480;
            {7'd40,7'd88}:		p = 14'd3520;
            {7'd40,7'd89}:		p = 14'd3560;
            {7'd40,7'd90}:		p = 14'd3600;
            {7'd40,7'd91}:		p = 14'd3640;
            {7'd40,7'd92}:		p = 14'd3680;
            {7'd40,7'd93}:		p = 14'd3720;
            {7'd40,7'd94}:		p = 14'd3760;
            {7'd40,7'd95}:		p = 14'd3800;
            {7'd40,7'd96}:		p = 14'd3840;
            {7'd40,7'd97}:		p = 14'd3880;
            {7'd40,7'd98}:		p = 14'd3920;
            {7'd40,7'd99}:		p = 14'd3960;
            {7'd40,7'd100}:		p = 14'd4000;
            {7'd40,7'd101}:		p = 14'd4040;
            {7'd40,7'd102}:		p = 14'd4080;
            {7'd40,7'd103}:		p = 14'd4120;
            {7'd40,7'd104}:		p = 14'd4160;
            {7'd40,7'd105}:		p = 14'd4200;
            {7'd40,7'd106}:		p = 14'd4240;
            {7'd40,7'd107}:		p = 14'd4280;
            {7'd40,7'd108}:		p = 14'd4320;
            {7'd40,7'd109}:		p = 14'd4360;
            {7'd40,7'd110}:		p = 14'd4400;
            {7'd40,7'd111}:		p = 14'd4440;
            {7'd40,7'd112}:		p = 14'd4480;
            {7'd40,7'd113}:		p = 14'd4520;
            {7'd40,7'd114}:		p = 14'd4560;
            {7'd40,7'd115}:		p = 14'd4600;
            {7'd40,7'd116}:		p = 14'd4640;
            {7'd40,7'd117}:		p = 14'd4680;
            {7'd40,7'd118}:		p = 14'd4720;
            {7'd40,7'd119}:		p = 14'd4760;
            {7'd40,7'd120}:		p = 14'd4800;
            {7'd40,7'd121}:		p = 14'd4840;
            {7'd40,7'd122}:		p = 14'd4880;
            {7'd40,7'd123}:		p = 14'd4920;
            {7'd40,7'd124}:		p = 14'd4960;
            {7'd40,7'd125}:		p = 14'd5000;
            {7'd40,7'd126}:		p = 14'd5040;
            {7'd40,7'd127}:		p = 14'd5080;
            {7'd41,7'd0}:		p = 14'd0;
            {7'd41,7'd1}:		p = 14'd41;
            {7'd41,7'd2}:		p = 14'd82;
            {7'd41,7'd3}:		p = 14'd123;
            {7'd41,7'd4}:		p = 14'd164;
            {7'd41,7'd5}:		p = 14'd205;
            {7'd41,7'd6}:		p = 14'd246;
            {7'd41,7'd7}:		p = 14'd287;
            {7'd41,7'd8}:		p = 14'd328;
            {7'd41,7'd9}:		p = 14'd369;
            {7'd41,7'd10}:		p = 14'd410;
            {7'd41,7'd11}:		p = 14'd451;
            {7'd41,7'd12}:		p = 14'd492;
            {7'd41,7'd13}:		p = 14'd533;
            {7'd41,7'd14}:		p = 14'd574;
            {7'd41,7'd15}:		p = 14'd615;
            {7'd41,7'd16}:		p = 14'd656;
            {7'd41,7'd17}:		p = 14'd697;
            {7'd41,7'd18}:		p = 14'd738;
            {7'd41,7'd19}:		p = 14'd779;
            {7'd41,7'd20}:		p = 14'd820;
            {7'd41,7'd21}:		p = 14'd861;
            {7'd41,7'd22}:		p = 14'd902;
            {7'd41,7'd23}:		p = 14'd943;
            {7'd41,7'd24}:		p = 14'd984;
            {7'd41,7'd25}:		p = 14'd1025;
            {7'd41,7'd26}:		p = 14'd1066;
            {7'd41,7'd27}:		p = 14'd1107;
            {7'd41,7'd28}:		p = 14'd1148;
            {7'd41,7'd29}:		p = 14'd1189;
            {7'd41,7'd30}:		p = 14'd1230;
            {7'd41,7'd31}:		p = 14'd1271;
            {7'd41,7'd32}:		p = 14'd1312;
            {7'd41,7'd33}:		p = 14'd1353;
            {7'd41,7'd34}:		p = 14'd1394;
            {7'd41,7'd35}:		p = 14'd1435;
            {7'd41,7'd36}:		p = 14'd1476;
            {7'd41,7'd37}:		p = 14'd1517;
            {7'd41,7'd38}:		p = 14'd1558;
            {7'd41,7'd39}:		p = 14'd1599;
            {7'd41,7'd40}:		p = 14'd1640;
            {7'd41,7'd41}:		p = 14'd1681;
            {7'd41,7'd42}:		p = 14'd1722;
            {7'd41,7'd43}:		p = 14'd1763;
            {7'd41,7'd44}:		p = 14'd1804;
            {7'd41,7'd45}:		p = 14'd1845;
            {7'd41,7'd46}:		p = 14'd1886;
            {7'd41,7'd47}:		p = 14'd1927;
            {7'd41,7'd48}:		p = 14'd1968;
            {7'd41,7'd49}:		p = 14'd2009;
            {7'd41,7'd50}:		p = 14'd2050;
            {7'd41,7'd51}:		p = 14'd2091;
            {7'd41,7'd52}:		p = 14'd2132;
            {7'd41,7'd53}:		p = 14'd2173;
            {7'd41,7'd54}:		p = 14'd2214;
            {7'd41,7'd55}:		p = 14'd2255;
            {7'd41,7'd56}:		p = 14'd2296;
            {7'd41,7'd57}:		p = 14'd2337;
            {7'd41,7'd58}:		p = 14'd2378;
            {7'd41,7'd59}:		p = 14'd2419;
            {7'd41,7'd60}:		p = 14'd2460;
            {7'd41,7'd61}:		p = 14'd2501;
            {7'd41,7'd62}:		p = 14'd2542;
            {7'd41,7'd63}:		p = 14'd2583;
            {7'd41,7'd64}:		p = 14'd2624;
            {7'd41,7'd65}:		p = 14'd2665;
            {7'd41,7'd66}:		p = 14'd2706;
            {7'd41,7'd67}:		p = 14'd2747;
            {7'd41,7'd68}:		p = 14'd2788;
            {7'd41,7'd69}:		p = 14'd2829;
            {7'd41,7'd70}:		p = 14'd2870;
            {7'd41,7'd71}:		p = 14'd2911;
            {7'd41,7'd72}:		p = 14'd2952;
            {7'd41,7'd73}:		p = 14'd2993;
            {7'd41,7'd74}:		p = 14'd3034;
            {7'd41,7'd75}:		p = 14'd3075;
            {7'd41,7'd76}:		p = 14'd3116;
            {7'd41,7'd77}:		p = 14'd3157;
            {7'd41,7'd78}:		p = 14'd3198;
            {7'd41,7'd79}:		p = 14'd3239;
            {7'd41,7'd80}:		p = 14'd3280;
            {7'd41,7'd81}:		p = 14'd3321;
            {7'd41,7'd82}:		p = 14'd3362;
            {7'd41,7'd83}:		p = 14'd3403;
            {7'd41,7'd84}:		p = 14'd3444;
            {7'd41,7'd85}:		p = 14'd3485;
            {7'd41,7'd86}:		p = 14'd3526;
            {7'd41,7'd87}:		p = 14'd3567;
            {7'd41,7'd88}:		p = 14'd3608;
            {7'd41,7'd89}:		p = 14'd3649;
            {7'd41,7'd90}:		p = 14'd3690;
            {7'd41,7'd91}:		p = 14'd3731;
            {7'd41,7'd92}:		p = 14'd3772;
            {7'd41,7'd93}:		p = 14'd3813;
            {7'd41,7'd94}:		p = 14'd3854;
            {7'd41,7'd95}:		p = 14'd3895;
            {7'd41,7'd96}:		p = 14'd3936;
            {7'd41,7'd97}:		p = 14'd3977;
            {7'd41,7'd98}:		p = 14'd4018;
            {7'd41,7'd99}:		p = 14'd4059;
            {7'd41,7'd100}:		p = 14'd4100;
            {7'd41,7'd101}:		p = 14'd4141;
            {7'd41,7'd102}:		p = 14'd4182;
            {7'd41,7'd103}:		p = 14'd4223;
            {7'd41,7'd104}:		p = 14'd4264;
            {7'd41,7'd105}:		p = 14'd4305;
            {7'd41,7'd106}:		p = 14'd4346;
            {7'd41,7'd107}:		p = 14'd4387;
            {7'd41,7'd108}:		p = 14'd4428;
            {7'd41,7'd109}:		p = 14'd4469;
            {7'd41,7'd110}:		p = 14'd4510;
            {7'd41,7'd111}:		p = 14'd4551;
            {7'd41,7'd112}:		p = 14'd4592;
            {7'd41,7'd113}:		p = 14'd4633;
            {7'd41,7'd114}:		p = 14'd4674;
            {7'd41,7'd115}:		p = 14'd4715;
            {7'd41,7'd116}:		p = 14'd4756;
            {7'd41,7'd117}:		p = 14'd4797;
            {7'd41,7'd118}:		p = 14'd4838;
            {7'd41,7'd119}:		p = 14'd4879;
            {7'd41,7'd120}:		p = 14'd4920;
            {7'd41,7'd121}:		p = 14'd4961;
            {7'd41,7'd122}:		p = 14'd5002;
            {7'd41,7'd123}:		p = 14'd5043;
            {7'd41,7'd124}:		p = 14'd5084;
            {7'd41,7'd125}:		p = 14'd5125;
            {7'd41,7'd126}:		p = 14'd5166;
            {7'd41,7'd127}:		p = 14'd5207;
            {7'd42,7'd0}:		p = 14'd0;
            {7'd42,7'd1}:		p = 14'd42;
            {7'd42,7'd2}:		p = 14'd84;
            {7'd42,7'd3}:		p = 14'd126;
            {7'd42,7'd4}:		p = 14'd168;
            {7'd42,7'd5}:		p = 14'd210;
            {7'd42,7'd6}:		p = 14'd252;
            {7'd42,7'd7}:		p = 14'd294;
            {7'd42,7'd8}:		p = 14'd336;
            {7'd42,7'd9}:		p = 14'd378;
            {7'd42,7'd10}:		p = 14'd420;
            {7'd42,7'd11}:		p = 14'd462;
            {7'd42,7'd12}:		p = 14'd504;
            {7'd42,7'd13}:		p = 14'd546;
            {7'd42,7'd14}:		p = 14'd588;
            {7'd42,7'd15}:		p = 14'd630;
            {7'd42,7'd16}:		p = 14'd672;
            {7'd42,7'd17}:		p = 14'd714;
            {7'd42,7'd18}:		p = 14'd756;
            {7'd42,7'd19}:		p = 14'd798;
            {7'd42,7'd20}:		p = 14'd840;
            {7'd42,7'd21}:		p = 14'd882;
            {7'd42,7'd22}:		p = 14'd924;
            {7'd42,7'd23}:		p = 14'd966;
            {7'd42,7'd24}:		p = 14'd1008;
            {7'd42,7'd25}:		p = 14'd1050;
            {7'd42,7'd26}:		p = 14'd1092;
            {7'd42,7'd27}:		p = 14'd1134;
            {7'd42,7'd28}:		p = 14'd1176;
            {7'd42,7'd29}:		p = 14'd1218;
            {7'd42,7'd30}:		p = 14'd1260;
            {7'd42,7'd31}:		p = 14'd1302;
            {7'd42,7'd32}:		p = 14'd1344;
            {7'd42,7'd33}:		p = 14'd1386;
            {7'd42,7'd34}:		p = 14'd1428;
            {7'd42,7'd35}:		p = 14'd1470;
            {7'd42,7'd36}:		p = 14'd1512;
            {7'd42,7'd37}:		p = 14'd1554;
            {7'd42,7'd38}:		p = 14'd1596;
            {7'd42,7'd39}:		p = 14'd1638;
            {7'd42,7'd40}:		p = 14'd1680;
            {7'd42,7'd41}:		p = 14'd1722;
            {7'd42,7'd42}:		p = 14'd1764;
            {7'd42,7'd43}:		p = 14'd1806;
            {7'd42,7'd44}:		p = 14'd1848;
            {7'd42,7'd45}:		p = 14'd1890;
            {7'd42,7'd46}:		p = 14'd1932;
            {7'd42,7'd47}:		p = 14'd1974;
            {7'd42,7'd48}:		p = 14'd2016;
            {7'd42,7'd49}:		p = 14'd2058;
            {7'd42,7'd50}:		p = 14'd2100;
            {7'd42,7'd51}:		p = 14'd2142;
            {7'd42,7'd52}:		p = 14'd2184;
            {7'd42,7'd53}:		p = 14'd2226;
            {7'd42,7'd54}:		p = 14'd2268;
            {7'd42,7'd55}:		p = 14'd2310;
            {7'd42,7'd56}:		p = 14'd2352;
            {7'd42,7'd57}:		p = 14'd2394;
            {7'd42,7'd58}:		p = 14'd2436;
            {7'd42,7'd59}:		p = 14'd2478;
            {7'd42,7'd60}:		p = 14'd2520;
            {7'd42,7'd61}:		p = 14'd2562;
            {7'd42,7'd62}:		p = 14'd2604;
            {7'd42,7'd63}:		p = 14'd2646;
            {7'd42,7'd64}:		p = 14'd2688;
            {7'd42,7'd65}:		p = 14'd2730;
            {7'd42,7'd66}:		p = 14'd2772;
            {7'd42,7'd67}:		p = 14'd2814;
            {7'd42,7'd68}:		p = 14'd2856;
            {7'd42,7'd69}:		p = 14'd2898;
            {7'd42,7'd70}:		p = 14'd2940;
            {7'd42,7'd71}:		p = 14'd2982;
            {7'd42,7'd72}:		p = 14'd3024;
            {7'd42,7'd73}:		p = 14'd3066;
            {7'd42,7'd74}:		p = 14'd3108;
            {7'd42,7'd75}:		p = 14'd3150;
            {7'd42,7'd76}:		p = 14'd3192;
            {7'd42,7'd77}:		p = 14'd3234;
            {7'd42,7'd78}:		p = 14'd3276;
            {7'd42,7'd79}:		p = 14'd3318;
            {7'd42,7'd80}:		p = 14'd3360;
            {7'd42,7'd81}:		p = 14'd3402;
            {7'd42,7'd82}:		p = 14'd3444;
            {7'd42,7'd83}:		p = 14'd3486;
            {7'd42,7'd84}:		p = 14'd3528;
            {7'd42,7'd85}:		p = 14'd3570;
            {7'd42,7'd86}:		p = 14'd3612;
            {7'd42,7'd87}:		p = 14'd3654;
            {7'd42,7'd88}:		p = 14'd3696;
            {7'd42,7'd89}:		p = 14'd3738;
            {7'd42,7'd90}:		p = 14'd3780;
            {7'd42,7'd91}:		p = 14'd3822;
            {7'd42,7'd92}:		p = 14'd3864;
            {7'd42,7'd93}:		p = 14'd3906;
            {7'd42,7'd94}:		p = 14'd3948;
            {7'd42,7'd95}:		p = 14'd3990;
            {7'd42,7'd96}:		p = 14'd4032;
            {7'd42,7'd97}:		p = 14'd4074;
            {7'd42,7'd98}:		p = 14'd4116;
            {7'd42,7'd99}:		p = 14'd4158;
            {7'd42,7'd100}:		p = 14'd4200;
            {7'd42,7'd101}:		p = 14'd4242;
            {7'd42,7'd102}:		p = 14'd4284;
            {7'd42,7'd103}:		p = 14'd4326;
            {7'd42,7'd104}:		p = 14'd4368;
            {7'd42,7'd105}:		p = 14'd4410;
            {7'd42,7'd106}:		p = 14'd4452;
            {7'd42,7'd107}:		p = 14'd4494;
            {7'd42,7'd108}:		p = 14'd4536;
            {7'd42,7'd109}:		p = 14'd4578;
            {7'd42,7'd110}:		p = 14'd4620;
            {7'd42,7'd111}:		p = 14'd4662;
            {7'd42,7'd112}:		p = 14'd4704;
            {7'd42,7'd113}:		p = 14'd4746;
            {7'd42,7'd114}:		p = 14'd4788;
            {7'd42,7'd115}:		p = 14'd4830;
            {7'd42,7'd116}:		p = 14'd4872;
            {7'd42,7'd117}:		p = 14'd4914;
            {7'd42,7'd118}:		p = 14'd4956;
            {7'd42,7'd119}:		p = 14'd4998;
            {7'd42,7'd120}:		p = 14'd5040;
            {7'd42,7'd121}:		p = 14'd5082;
            {7'd42,7'd122}:		p = 14'd5124;
            {7'd42,7'd123}:		p = 14'd5166;
            {7'd42,7'd124}:		p = 14'd5208;
            {7'd42,7'd125}:		p = 14'd5250;
            {7'd42,7'd126}:		p = 14'd5292;
            {7'd42,7'd127}:		p = 14'd5334;
            {7'd43,7'd0}:		p = 14'd0;
            {7'd43,7'd1}:		p = 14'd43;
            {7'd43,7'd2}:		p = 14'd86;
            {7'd43,7'd3}:		p = 14'd129;
            {7'd43,7'd4}:		p = 14'd172;
            {7'd43,7'd5}:		p = 14'd215;
            {7'd43,7'd6}:		p = 14'd258;
            {7'd43,7'd7}:		p = 14'd301;
            {7'd43,7'd8}:		p = 14'd344;
            {7'd43,7'd9}:		p = 14'd387;
            {7'd43,7'd10}:		p = 14'd430;
            {7'd43,7'd11}:		p = 14'd473;
            {7'd43,7'd12}:		p = 14'd516;
            {7'd43,7'd13}:		p = 14'd559;
            {7'd43,7'd14}:		p = 14'd602;
            {7'd43,7'd15}:		p = 14'd645;
            {7'd43,7'd16}:		p = 14'd688;
            {7'd43,7'd17}:		p = 14'd731;
            {7'd43,7'd18}:		p = 14'd774;
            {7'd43,7'd19}:		p = 14'd817;
            {7'd43,7'd20}:		p = 14'd860;
            {7'd43,7'd21}:		p = 14'd903;
            {7'd43,7'd22}:		p = 14'd946;
            {7'd43,7'd23}:		p = 14'd989;
            {7'd43,7'd24}:		p = 14'd1032;
            {7'd43,7'd25}:		p = 14'd1075;
            {7'd43,7'd26}:		p = 14'd1118;
            {7'd43,7'd27}:		p = 14'd1161;
            {7'd43,7'd28}:		p = 14'd1204;
            {7'd43,7'd29}:		p = 14'd1247;
            {7'd43,7'd30}:		p = 14'd1290;
            {7'd43,7'd31}:		p = 14'd1333;
            {7'd43,7'd32}:		p = 14'd1376;
            {7'd43,7'd33}:		p = 14'd1419;
            {7'd43,7'd34}:		p = 14'd1462;
            {7'd43,7'd35}:		p = 14'd1505;
            {7'd43,7'd36}:		p = 14'd1548;
            {7'd43,7'd37}:		p = 14'd1591;
            {7'd43,7'd38}:		p = 14'd1634;
            {7'd43,7'd39}:		p = 14'd1677;
            {7'd43,7'd40}:		p = 14'd1720;
            {7'd43,7'd41}:		p = 14'd1763;
            {7'd43,7'd42}:		p = 14'd1806;
            {7'd43,7'd43}:		p = 14'd1849;
            {7'd43,7'd44}:		p = 14'd1892;
            {7'd43,7'd45}:		p = 14'd1935;
            {7'd43,7'd46}:		p = 14'd1978;
            {7'd43,7'd47}:		p = 14'd2021;
            {7'd43,7'd48}:		p = 14'd2064;
            {7'd43,7'd49}:		p = 14'd2107;
            {7'd43,7'd50}:		p = 14'd2150;
            {7'd43,7'd51}:		p = 14'd2193;
            {7'd43,7'd52}:		p = 14'd2236;
            {7'd43,7'd53}:		p = 14'd2279;
            {7'd43,7'd54}:		p = 14'd2322;
            {7'd43,7'd55}:		p = 14'd2365;
            {7'd43,7'd56}:		p = 14'd2408;
            {7'd43,7'd57}:		p = 14'd2451;
            {7'd43,7'd58}:		p = 14'd2494;
            {7'd43,7'd59}:		p = 14'd2537;
            {7'd43,7'd60}:		p = 14'd2580;
            {7'd43,7'd61}:		p = 14'd2623;
            {7'd43,7'd62}:		p = 14'd2666;
            {7'd43,7'd63}:		p = 14'd2709;
            {7'd43,7'd64}:		p = 14'd2752;
            {7'd43,7'd65}:		p = 14'd2795;
            {7'd43,7'd66}:		p = 14'd2838;
            {7'd43,7'd67}:		p = 14'd2881;
            {7'd43,7'd68}:		p = 14'd2924;
            {7'd43,7'd69}:		p = 14'd2967;
            {7'd43,7'd70}:		p = 14'd3010;
            {7'd43,7'd71}:		p = 14'd3053;
            {7'd43,7'd72}:		p = 14'd3096;
            {7'd43,7'd73}:		p = 14'd3139;
            {7'd43,7'd74}:		p = 14'd3182;
            {7'd43,7'd75}:		p = 14'd3225;
            {7'd43,7'd76}:		p = 14'd3268;
            {7'd43,7'd77}:		p = 14'd3311;
            {7'd43,7'd78}:		p = 14'd3354;
            {7'd43,7'd79}:		p = 14'd3397;
            {7'd43,7'd80}:		p = 14'd3440;
            {7'd43,7'd81}:		p = 14'd3483;
            {7'd43,7'd82}:		p = 14'd3526;
            {7'd43,7'd83}:		p = 14'd3569;
            {7'd43,7'd84}:		p = 14'd3612;
            {7'd43,7'd85}:		p = 14'd3655;
            {7'd43,7'd86}:		p = 14'd3698;
            {7'd43,7'd87}:		p = 14'd3741;
            {7'd43,7'd88}:		p = 14'd3784;
            {7'd43,7'd89}:		p = 14'd3827;
            {7'd43,7'd90}:		p = 14'd3870;
            {7'd43,7'd91}:		p = 14'd3913;
            {7'd43,7'd92}:		p = 14'd3956;
            {7'd43,7'd93}:		p = 14'd3999;
            {7'd43,7'd94}:		p = 14'd4042;
            {7'd43,7'd95}:		p = 14'd4085;
            {7'd43,7'd96}:		p = 14'd4128;
            {7'd43,7'd97}:		p = 14'd4171;
            {7'd43,7'd98}:		p = 14'd4214;
            {7'd43,7'd99}:		p = 14'd4257;
            {7'd43,7'd100}:		p = 14'd4300;
            {7'd43,7'd101}:		p = 14'd4343;
            {7'd43,7'd102}:		p = 14'd4386;
            {7'd43,7'd103}:		p = 14'd4429;
            {7'd43,7'd104}:		p = 14'd4472;
            {7'd43,7'd105}:		p = 14'd4515;
            {7'd43,7'd106}:		p = 14'd4558;
            {7'd43,7'd107}:		p = 14'd4601;
            {7'd43,7'd108}:		p = 14'd4644;
            {7'd43,7'd109}:		p = 14'd4687;
            {7'd43,7'd110}:		p = 14'd4730;
            {7'd43,7'd111}:		p = 14'd4773;
            {7'd43,7'd112}:		p = 14'd4816;
            {7'd43,7'd113}:		p = 14'd4859;
            {7'd43,7'd114}:		p = 14'd4902;
            {7'd43,7'd115}:		p = 14'd4945;
            {7'd43,7'd116}:		p = 14'd4988;
            {7'd43,7'd117}:		p = 14'd5031;
            {7'd43,7'd118}:		p = 14'd5074;
            {7'd43,7'd119}:		p = 14'd5117;
            {7'd43,7'd120}:		p = 14'd5160;
            {7'd43,7'd121}:		p = 14'd5203;
            {7'd43,7'd122}:		p = 14'd5246;
            {7'd43,7'd123}:		p = 14'd5289;
            {7'd43,7'd124}:		p = 14'd5332;
            {7'd43,7'd125}:		p = 14'd5375;
            {7'd43,7'd126}:		p = 14'd5418;
            {7'd43,7'd127}:		p = 14'd5461;
            {7'd44,7'd0}:		p = 14'd0;
            {7'd44,7'd1}:		p = 14'd44;
            {7'd44,7'd2}:		p = 14'd88;
            {7'd44,7'd3}:		p = 14'd132;
            {7'd44,7'd4}:		p = 14'd176;
            {7'd44,7'd5}:		p = 14'd220;
            {7'd44,7'd6}:		p = 14'd264;
            {7'd44,7'd7}:		p = 14'd308;
            {7'd44,7'd8}:		p = 14'd352;
            {7'd44,7'd9}:		p = 14'd396;
            {7'd44,7'd10}:		p = 14'd440;
            {7'd44,7'd11}:		p = 14'd484;
            {7'd44,7'd12}:		p = 14'd528;
            {7'd44,7'd13}:		p = 14'd572;
            {7'd44,7'd14}:		p = 14'd616;
            {7'd44,7'd15}:		p = 14'd660;
            {7'd44,7'd16}:		p = 14'd704;
            {7'd44,7'd17}:		p = 14'd748;
            {7'd44,7'd18}:		p = 14'd792;
            {7'd44,7'd19}:		p = 14'd836;
            {7'd44,7'd20}:		p = 14'd880;
            {7'd44,7'd21}:		p = 14'd924;
            {7'd44,7'd22}:		p = 14'd968;
            {7'd44,7'd23}:		p = 14'd1012;
            {7'd44,7'd24}:		p = 14'd1056;
            {7'd44,7'd25}:		p = 14'd1100;
            {7'd44,7'd26}:		p = 14'd1144;
            {7'd44,7'd27}:		p = 14'd1188;
            {7'd44,7'd28}:		p = 14'd1232;
            {7'd44,7'd29}:		p = 14'd1276;
            {7'd44,7'd30}:		p = 14'd1320;
            {7'd44,7'd31}:		p = 14'd1364;
            {7'd44,7'd32}:		p = 14'd1408;
            {7'd44,7'd33}:		p = 14'd1452;
            {7'd44,7'd34}:		p = 14'd1496;
            {7'd44,7'd35}:		p = 14'd1540;
            {7'd44,7'd36}:		p = 14'd1584;
            {7'd44,7'd37}:		p = 14'd1628;
            {7'd44,7'd38}:		p = 14'd1672;
            {7'd44,7'd39}:		p = 14'd1716;
            {7'd44,7'd40}:		p = 14'd1760;
            {7'd44,7'd41}:		p = 14'd1804;
            {7'd44,7'd42}:		p = 14'd1848;
            {7'd44,7'd43}:		p = 14'd1892;
            {7'd44,7'd44}:		p = 14'd1936;
            {7'd44,7'd45}:		p = 14'd1980;
            {7'd44,7'd46}:		p = 14'd2024;
            {7'd44,7'd47}:		p = 14'd2068;
            {7'd44,7'd48}:		p = 14'd2112;
            {7'd44,7'd49}:		p = 14'd2156;
            {7'd44,7'd50}:		p = 14'd2200;
            {7'd44,7'd51}:		p = 14'd2244;
            {7'd44,7'd52}:		p = 14'd2288;
            {7'd44,7'd53}:		p = 14'd2332;
            {7'd44,7'd54}:		p = 14'd2376;
            {7'd44,7'd55}:		p = 14'd2420;
            {7'd44,7'd56}:		p = 14'd2464;
            {7'd44,7'd57}:		p = 14'd2508;
            {7'd44,7'd58}:		p = 14'd2552;
            {7'd44,7'd59}:		p = 14'd2596;
            {7'd44,7'd60}:		p = 14'd2640;
            {7'd44,7'd61}:		p = 14'd2684;
            {7'd44,7'd62}:		p = 14'd2728;
            {7'd44,7'd63}:		p = 14'd2772;
            {7'd44,7'd64}:		p = 14'd2816;
            {7'd44,7'd65}:		p = 14'd2860;
            {7'd44,7'd66}:		p = 14'd2904;
            {7'd44,7'd67}:		p = 14'd2948;
            {7'd44,7'd68}:		p = 14'd2992;
            {7'd44,7'd69}:		p = 14'd3036;
            {7'd44,7'd70}:		p = 14'd3080;
            {7'd44,7'd71}:		p = 14'd3124;
            {7'd44,7'd72}:		p = 14'd3168;
            {7'd44,7'd73}:		p = 14'd3212;
            {7'd44,7'd74}:		p = 14'd3256;
            {7'd44,7'd75}:		p = 14'd3300;
            {7'd44,7'd76}:		p = 14'd3344;
            {7'd44,7'd77}:		p = 14'd3388;
            {7'd44,7'd78}:		p = 14'd3432;
            {7'd44,7'd79}:		p = 14'd3476;
            {7'd44,7'd80}:		p = 14'd3520;
            {7'd44,7'd81}:		p = 14'd3564;
            {7'd44,7'd82}:		p = 14'd3608;
            {7'd44,7'd83}:		p = 14'd3652;
            {7'd44,7'd84}:		p = 14'd3696;
            {7'd44,7'd85}:		p = 14'd3740;
            {7'd44,7'd86}:		p = 14'd3784;
            {7'd44,7'd87}:		p = 14'd3828;
            {7'd44,7'd88}:		p = 14'd3872;
            {7'd44,7'd89}:		p = 14'd3916;
            {7'd44,7'd90}:		p = 14'd3960;
            {7'd44,7'd91}:		p = 14'd4004;
            {7'd44,7'd92}:		p = 14'd4048;
            {7'd44,7'd93}:		p = 14'd4092;
            {7'd44,7'd94}:		p = 14'd4136;
            {7'd44,7'd95}:		p = 14'd4180;
            {7'd44,7'd96}:		p = 14'd4224;
            {7'd44,7'd97}:		p = 14'd4268;
            {7'd44,7'd98}:		p = 14'd4312;
            {7'd44,7'd99}:		p = 14'd4356;
            {7'd44,7'd100}:		p = 14'd4400;
            {7'd44,7'd101}:		p = 14'd4444;
            {7'd44,7'd102}:		p = 14'd4488;
            {7'd44,7'd103}:		p = 14'd4532;
            {7'd44,7'd104}:		p = 14'd4576;
            {7'd44,7'd105}:		p = 14'd4620;
            {7'd44,7'd106}:		p = 14'd4664;
            {7'd44,7'd107}:		p = 14'd4708;
            {7'd44,7'd108}:		p = 14'd4752;
            {7'd44,7'd109}:		p = 14'd4796;
            {7'd44,7'd110}:		p = 14'd4840;
            {7'd44,7'd111}:		p = 14'd4884;
            {7'd44,7'd112}:		p = 14'd4928;
            {7'd44,7'd113}:		p = 14'd4972;
            {7'd44,7'd114}:		p = 14'd5016;
            {7'd44,7'd115}:		p = 14'd5060;
            {7'd44,7'd116}:		p = 14'd5104;
            {7'd44,7'd117}:		p = 14'd5148;
            {7'd44,7'd118}:		p = 14'd5192;
            {7'd44,7'd119}:		p = 14'd5236;
            {7'd44,7'd120}:		p = 14'd5280;
            {7'd44,7'd121}:		p = 14'd5324;
            {7'd44,7'd122}:		p = 14'd5368;
            {7'd44,7'd123}:		p = 14'd5412;
            {7'd44,7'd124}:		p = 14'd5456;
            {7'd44,7'd125}:		p = 14'd5500;
            {7'd44,7'd126}:		p = 14'd5544;
            {7'd44,7'd127}:		p = 14'd5588;
            {7'd45,7'd0}:		p = 14'd0;
            {7'd45,7'd1}:		p = 14'd45;
            {7'd45,7'd2}:		p = 14'd90;
            {7'd45,7'd3}:		p = 14'd135;
            {7'd45,7'd4}:		p = 14'd180;
            {7'd45,7'd5}:		p = 14'd225;
            {7'd45,7'd6}:		p = 14'd270;
            {7'd45,7'd7}:		p = 14'd315;
            {7'd45,7'd8}:		p = 14'd360;
            {7'd45,7'd9}:		p = 14'd405;
            {7'd45,7'd10}:		p = 14'd450;
            {7'd45,7'd11}:		p = 14'd495;
            {7'd45,7'd12}:		p = 14'd540;
            {7'd45,7'd13}:		p = 14'd585;
            {7'd45,7'd14}:		p = 14'd630;
            {7'd45,7'd15}:		p = 14'd675;
            {7'd45,7'd16}:		p = 14'd720;
            {7'd45,7'd17}:		p = 14'd765;
            {7'd45,7'd18}:		p = 14'd810;
            {7'd45,7'd19}:		p = 14'd855;
            {7'd45,7'd20}:		p = 14'd900;
            {7'd45,7'd21}:		p = 14'd945;
            {7'd45,7'd22}:		p = 14'd990;
            {7'd45,7'd23}:		p = 14'd1035;
            {7'd45,7'd24}:		p = 14'd1080;
            {7'd45,7'd25}:		p = 14'd1125;
            {7'd45,7'd26}:		p = 14'd1170;
            {7'd45,7'd27}:		p = 14'd1215;
            {7'd45,7'd28}:		p = 14'd1260;
            {7'd45,7'd29}:		p = 14'd1305;
            {7'd45,7'd30}:		p = 14'd1350;
            {7'd45,7'd31}:		p = 14'd1395;
            {7'd45,7'd32}:		p = 14'd1440;
            {7'd45,7'd33}:		p = 14'd1485;
            {7'd45,7'd34}:		p = 14'd1530;
            {7'd45,7'd35}:		p = 14'd1575;
            {7'd45,7'd36}:		p = 14'd1620;
            {7'd45,7'd37}:		p = 14'd1665;
            {7'd45,7'd38}:		p = 14'd1710;
            {7'd45,7'd39}:		p = 14'd1755;
            {7'd45,7'd40}:		p = 14'd1800;
            {7'd45,7'd41}:		p = 14'd1845;
            {7'd45,7'd42}:		p = 14'd1890;
            {7'd45,7'd43}:		p = 14'd1935;
            {7'd45,7'd44}:		p = 14'd1980;
            {7'd45,7'd45}:		p = 14'd2025;
            {7'd45,7'd46}:		p = 14'd2070;
            {7'd45,7'd47}:		p = 14'd2115;
            {7'd45,7'd48}:		p = 14'd2160;
            {7'd45,7'd49}:		p = 14'd2205;
            {7'd45,7'd50}:		p = 14'd2250;
            {7'd45,7'd51}:		p = 14'd2295;
            {7'd45,7'd52}:		p = 14'd2340;
            {7'd45,7'd53}:		p = 14'd2385;
            {7'd45,7'd54}:		p = 14'd2430;
            {7'd45,7'd55}:		p = 14'd2475;
            {7'd45,7'd56}:		p = 14'd2520;
            {7'd45,7'd57}:		p = 14'd2565;
            {7'd45,7'd58}:		p = 14'd2610;
            {7'd45,7'd59}:		p = 14'd2655;
            {7'd45,7'd60}:		p = 14'd2700;
            {7'd45,7'd61}:		p = 14'd2745;
            {7'd45,7'd62}:		p = 14'd2790;
            {7'd45,7'd63}:		p = 14'd2835;
            {7'd45,7'd64}:		p = 14'd2880;
            {7'd45,7'd65}:		p = 14'd2925;
            {7'd45,7'd66}:		p = 14'd2970;
            {7'd45,7'd67}:		p = 14'd3015;
            {7'd45,7'd68}:		p = 14'd3060;
            {7'd45,7'd69}:		p = 14'd3105;
            {7'd45,7'd70}:		p = 14'd3150;
            {7'd45,7'd71}:		p = 14'd3195;
            {7'd45,7'd72}:		p = 14'd3240;
            {7'd45,7'd73}:		p = 14'd3285;
            {7'd45,7'd74}:		p = 14'd3330;
            {7'd45,7'd75}:		p = 14'd3375;
            {7'd45,7'd76}:		p = 14'd3420;
            {7'd45,7'd77}:		p = 14'd3465;
            {7'd45,7'd78}:		p = 14'd3510;
            {7'd45,7'd79}:		p = 14'd3555;
            {7'd45,7'd80}:		p = 14'd3600;
            {7'd45,7'd81}:		p = 14'd3645;
            {7'd45,7'd82}:		p = 14'd3690;
            {7'd45,7'd83}:		p = 14'd3735;
            {7'd45,7'd84}:		p = 14'd3780;
            {7'd45,7'd85}:		p = 14'd3825;
            {7'd45,7'd86}:		p = 14'd3870;
            {7'd45,7'd87}:		p = 14'd3915;
            {7'd45,7'd88}:		p = 14'd3960;
            {7'd45,7'd89}:		p = 14'd4005;
            {7'd45,7'd90}:		p = 14'd4050;
            {7'd45,7'd91}:		p = 14'd4095;
            {7'd45,7'd92}:		p = 14'd4140;
            {7'd45,7'd93}:		p = 14'd4185;
            {7'd45,7'd94}:		p = 14'd4230;
            {7'd45,7'd95}:		p = 14'd4275;
            {7'd45,7'd96}:		p = 14'd4320;
            {7'd45,7'd97}:		p = 14'd4365;
            {7'd45,7'd98}:		p = 14'd4410;
            {7'd45,7'd99}:		p = 14'd4455;
            {7'd45,7'd100}:		p = 14'd4500;
            {7'd45,7'd101}:		p = 14'd4545;
            {7'd45,7'd102}:		p = 14'd4590;
            {7'd45,7'd103}:		p = 14'd4635;
            {7'd45,7'd104}:		p = 14'd4680;
            {7'd45,7'd105}:		p = 14'd4725;
            {7'd45,7'd106}:		p = 14'd4770;
            {7'd45,7'd107}:		p = 14'd4815;
            {7'd45,7'd108}:		p = 14'd4860;
            {7'd45,7'd109}:		p = 14'd4905;
            {7'd45,7'd110}:		p = 14'd4950;
            {7'd45,7'd111}:		p = 14'd4995;
            {7'd45,7'd112}:		p = 14'd5040;
            {7'd45,7'd113}:		p = 14'd5085;
            {7'd45,7'd114}:		p = 14'd5130;
            {7'd45,7'd115}:		p = 14'd5175;
            {7'd45,7'd116}:		p = 14'd5220;
            {7'd45,7'd117}:		p = 14'd5265;
            {7'd45,7'd118}:		p = 14'd5310;
            {7'd45,7'd119}:		p = 14'd5355;
            {7'd45,7'd120}:		p = 14'd5400;
            {7'd45,7'd121}:		p = 14'd5445;
            {7'd45,7'd122}:		p = 14'd5490;
            {7'd45,7'd123}:		p = 14'd5535;
            {7'd45,7'd124}:		p = 14'd5580;
            {7'd45,7'd125}:		p = 14'd5625;
            {7'd45,7'd126}:		p = 14'd5670;
            {7'd45,7'd127}:		p = 14'd5715;
            {7'd46,7'd0}:		p = 14'd0;
            {7'd46,7'd1}:		p = 14'd46;
            {7'd46,7'd2}:		p = 14'd92;
            {7'd46,7'd3}:		p = 14'd138;
            {7'd46,7'd4}:		p = 14'd184;
            {7'd46,7'd5}:		p = 14'd230;
            {7'd46,7'd6}:		p = 14'd276;
            {7'd46,7'd7}:		p = 14'd322;
            {7'd46,7'd8}:		p = 14'd368;
            {7'd46,7'd9}:		p = 14'd414;
            {7'd46,7'd10}:		p = 14'd460;
            {7'd46,7'd11}:		p = 14'd506;
            {7'd46,7'd12}:		p = 14'd552;
            {7'd46,7'd13}:		p = 14'd598;
            {7'd46,7'd14}:		p = 14'd644;
            {7'd46,7'd15}:		p = 14'd690;
            {7'd46,7'd16}:		p = 14'd736;
            {7'd46,7'd17}:		p = 14'd782;
            {7'd46,7'd18}:		p = 14'd828;
            {7'd46,7'd19}:		p = 14'd874;
            {7'd46,7'd20}:		p = 14'd920;
            {7'd46,7'd21}:		p = 14'd966;
            {7'd46,7'd22}:		p = 14'd1012;
            {7'd46,7'd23}:		p = 14'd1058;
            {7'd46,7'd24}:		p = 14'd1104;
            {7'd46,7'd25}:		p = 14'd1150;
            {7'd46,7'd26}:		p = 14'd1196;
            {7'd46,7'd27}:		p = 14'd1242;
            {7'd46,7'd28}:		p = 14'd1288;
            {7'd46,7'd29}:		p = 14'd1334;
            {7'd46,7'd30}:		p = 14'd1380;
            {7'd46,7'd31}:		p = 14'd1426;
            {7'd46,7'd32}:		p = 14'd1472;
            {7'd46,7'd33}:		p = 14'd1518;
            {7'd46,7'd34}:		p = 14'd1564;
            {7'd46,7'd35}:		p = 14'd1610;
            {7'd46,7'd36}:		p = 14'd1656;
            {7'd46,7'd37}:		p = 14'd1702;
            {7'd46,7'd38}:		p = 14'd1748;
            {7'd46,7'd39}:		p = 14'd1794;
            {7'd46,7'd40}:		p = 14'd1840;
            {7'd46,7'd41}:		p = 14'd1886;
            {7'd46,7'd42}:		p = 14'd1932;
            {7'd46,7'd43}:		p = 14'd1978;
            {7'd46,7'd44}:		p = 14'd2024;
            {7'd46,7'd45}:		p = 14'd2070;
            {7'd46,7'd46}:		p = 14'd2116;
            {7'd46,7'd47}:		p = 14'd2162;
            {7'd46,7'd48}:		p = 14'd2208;
            {7'd46,7'd49}:		p = 14'd2254;
            {7'd46,7'd50}:		p = 14'd2300;
            {7'd46,7'd51}:		p = 14'd2346;
            {7'd46,7'd52}:		p = 14'd2392;
            {7'd46,7'd53}:		p = 14'd2438;
            {7'd46,7'd54}:		p = 14'd2484;
            {7'd46,7'd55}:		p = 14'd2530;
            {7'd46,7'd56}:		p = 14'd2576;
            {7'd46,7'd57}:		p = 14'd2622;
            {7'd46,7'd58}:		p = 14'd2668;
            {7'd46,7'd59}:		p = 14'd2714;
            {7'd46,7'd60}:		p = 14'd2760;
            {7'd46,7'd61}:		p = 14'd2806;
            {7'd46,7'd62}:		p = 14'd2852;
            {7'd46,7'd63}:		p = 14'd2898;
            {7'd46,7'd64}:		p = 14'd2944;
            {7'd46,7'd65}:		p = 14'd2990;
            {7'd46,7'd66}:		p = 14'd3036;
            {7'd46,7'd67}:		p = 14'd3082;
            {7'd46,7'd68}:		p = 14'd3128;
            {7'd46,7'd69}:		p = 14'd3174;
            {7'd46,7'd70}:		p = 14'd3220;
            {7'd46,7'd71}:		p = 14'd3266;
            {7'd46,7'd72}:		p = 14'd3312;
            {7'd46,7'd73}:		p = 14'd3358;
            {7'd46,7'd74}:		p = 14'd3404;
            {7'd46,7'd75}:		p = 14'd3450;
            {7'd46,7'd76}:		p = 14'd3496;
            {7'd46,7'd77}:		p = 14'd3542;
            {7'd46,7'd78}:		p = 14'd3588;
            {7'd46,7'd79}:		p = 14'd3634;
            {7'd46,7'd80}:		p = 14'd3680;
            {7'd46,7'd81}:		p = 14'd3726;
            {7'd46,7'd82}:		p = 14'd3772;
            {7'd46,7'd83}:		p = 14'd3818;
            {7'd46,7'd84}:		p = 14'd3864;
            {7'd46,7'd85}:		p = 14'd3910;
            {7'd46,7'd86}:		p = 14'd3956;
            {7'd46,7'd87}:		p = 14'd4002;
            {7'd46,7'd88}:		p = 14'd4048;
            {7'd46,7'd89}:		p = 14'd4094;
            {7'd46,7'd90}:		p = 14'd4140;
            {7'd46,7'd91}:		p = 14'd4186;
            {7'd46,7'd92}:		p = 14'd4232;
            {7'd46,7'd93}:		p = 14'd4278;
            {7'd46,7'd94}:		p = 14'd4324;
            {7'd46,7'd95}:		p = 14'd4370;
            {7'd46,7'd96}:		p = 14'd4416;
            {7'd46,7'd97}:		p = 14'd4462;
            {7'd46,7'd98}:		p = 14'd4508;
            {7'd46,7'd99}:		p = 14'd4554;
            {7'd46,7'd100}:		p = 14'd4600;
            {7'd46,7'd101}:		p = 14'd4646;
            {7'd46,7'd102}:		p = 14'd4692;
            {7'd46,7'd103}:		p = 14'd4738;
            {7'd46,7'd104}:		p = 14'd4784;
            {7'd46,7'd105}:		p = 14'd4830;
            {7'd46,7'd106}:		p = 14'd4876;
            {7'd46,7'd107}:		p = 14'd4922;
            {7'd46,7'd108}:		p = 14'd4968;
            {7'd46,7'd109}:		p = 14'd5014;
            {7'd46,7'd110}:		p = 14'd5060;
            {7'd46,7'd111}:		p = 14'd5106;
            {7'd46,7'd112}:		p = 14'd5152;
            {7'd46,7'd113}:		p = 14'd5198;
            {7'd46,7'd114}:		p = 14'd5244;
            {7'd46,7'd115}:		p = 14'd5290;
            {7'd46,7'd116}:		p = 14'd5336;
            {7'd46,7'd117}:		p = 14'd5382;
            {7'd46,7'd118}:		p = 14'd5428;
            {7'd46,7'd119}:		p = 14'd5474;
            {7'd46,7'd120}:		p = 14'd5520;
            {7'd46,7'd121}:		p = 14'd5566;
            {7'd46,7'd122}:		p = 14'd5612;
            {7'd46,7'd123}:		p = 14'd5658;
            {7'd46,7'd124}:		p = 14'd5704;
            {7'd46,7'd125}:		p = 14'd5750;
            {7'd46,7'd126}:		p = 14'd5796;
            {7'd46,7'd127}:		p = 14'd5842;
            {7'd47,7'd0}:		p = 14'd0;
            {7'd47,7'd1}:		p = 14'd47;
            {7'd47,7'd2}:		p = 14'd94;
            {7'd47,7'd3}:		p = 14'd141;
            {7'd47,7'd4}:		p = 14'd188;
            {7'd47,7'd5}:		p = 14'd235;
            {7'd47,7'd6}:		p = 14'd282;
            {7'd47,7'd7}:		p = 14'd329;
            {7'd47,7'd8}:		p = 14'd376;
            {7'd47,7'd9}:		p = 14'd423;
            {7'd47,7'd10}:		p = 14'd470;
            {7'd47,7'd11}:		p = 14'd517;
            {7'd47,7'd12}:		p = 14'd564;
            {7'd47,7'd13}:		p = 14'd611;
            {7'd47,7'd14}:		p = 14'd658;
            {7'd47,7'd15}:		p = 14'd705;
            {7'd47,7'd16}:		p = 14'd752;
            {7'd47,7'd17}:		p = 14'd799;
            {7'd47,7'd18}:		p = 14'd846;
            {7'd47,7'd19}:		p = 14'd893;
            {7'd47,7'd20}:		p = 14'd940;
            {7'd47,7'd21}:		p = 14'd987;
            {7'd47,7'd22}:		p = 14'd1034;
            {7'd47,7'd23}:		p = 14'd1081;
            {7'd47,7'd24}:		p = 14'd1128;
            {7'd47,7'd25}:		p = 14'd1175;
            {7'd47,7'd26}:		p = 14'd1222;
            {7'd47,7'd27}:		p = 14'd1269;
            {7'd47,7'd28}:		p = 14'd1316;
            {7'd47,7'd29}:		p = 14'd1363;
            {7'd47,7'd30}:		p = 14'd1410;
            {7'd47,7'd31}:		p = 14'd1457;
            {7'd47,7'd32}:		p = 14'd1504;
            {7'd47,7'd33}:		p = 14'd1551;
            {7'd47,7'd34}:		p = 14'd1598;
            {7'd47,7'd35}:		p = 14'd1645;
            {7'd47,7'd36}:		p = 14'd1692;
            {7'd47,7'd37}:		p = 14'd1739;
            {7'd47,7'd38}:		p = 14'd1786;
            {7'd47,7'd39}:		p = 14'd1833;
            {7'd47,7'd40}:		p = 14'd1880;
            {7'd47,7'd41}:		p = 14'd1927;
            {7'd47,7'd42}:		p = 14'd1974;
            {7'd47,7'd43}:		p = 14'd2021;
            {7'd47,7'd44}:		p = 14'd2068;
            {7'd47,7'd45}:		p = 14'd2115;
            {7'd47,7'd46}:		p = 14'd2162;
            {7'd47,7'd47}:		p = 14'd2209;
            {7'd47,7'd48}:		p = 14'd2256;
            {7'd47,7'd49}:		p = 14'd2303;
            {7'd47,7'd50}:		p = 14'd2350;
            {7'd47,7'd51}:		p = 14'd2397;
            {7'd47,7'd52}:		p = 14'd2444;
            {7'd47,7'd53}:		p = 14'd2491;
            {7'd47,7'd54}:		p = 14'd2538;
            {7'd47,7'd55}:		p = 14'd2585;
            {7'd47,7'd56}:		p = 14'd2632;
            {7'd47,7'd57}:		p = 14'd2679;
            {7'd47,7'd58}:		p = 14'd2726;
            {7'd47,7'd59}:		p = 14'd2773;
            {7'd47,7'd60}:		p = 14'd2820;
            {7'd47,7'd61}:		p = 14'd2867;
            {7'd47,7'd62}:		p = 14'd2914;
            {7'd47,7'd63}:		p = 14'd2961;
            {7'd47,7'd64}:		p = 14'd3008;
            {7'd47,7'd65}:		p = 14'd3055;
            {7'd47,7'd66}:		p = 14'd3102;
            {7'd47,7'd67}:		p = 14'd3149;
            {7'd47,7'd68}:		p = 14'd3196;
            {7'd47,7'd69}:		p = 14'd3243;
            {7'd47,7'd70}:		p = 14'd3290;
            {7'd47,7'd71}:		p = 14'd3337;
            {7'd47,7'd72}:		p = 14'd3384;
            {7'd47,7'd73}:		p = 14'd3431;
            {7'd47,7'd74}:		p = 14'd3478;
            {7'd47,7'd75}:		p = 14'd3525;
            {7'd47,7'd76}:		p = 14'd3572;
            {7'd47,7'd77}:		p = 14'd3619;
            {7'd47,7'd78}:		p = 14'd3666;
            {7'd47,7'd79}:		p = 14'd3713;
            {7'd47,7'd80}:		p = 14'd3760;
            {7'd47,7'd81}:		p = 14'd3807;
            {7'd47,7'd82}:		p = 14'd3854;
            {7'd47,7'd83}:		p = 14'd3901;
            {7'd47,7'd84}:		p = 14'd3948;
            {7'd47,7'd85}:		p = 14'd3995;
            {7'd47,7'd86}:		p = 14'd4042;
            {7'd47,7'd87}:		p = 14'd4089;
            {7'd47,7'd88}:		p = 14'd4136;
            {7'd47,7'd89}:		p = 14'd4183;
            {7'd47,7'd90}:		p = 14'd4230;
            {7'd47,7'd91}:		p = 14'd4277;
            {7'd47,7'd92}:		p = 14'd4324;
            {7'd47,7'd93}:		p = 14'd4371;
            {7'd47,7'd94}:		p = 14'd4418;
            {7'd47,7'd95}:		p = 14'd4465;
            {7'd47,7'd96}:		p = 14'd4512;
            {7'd47,7'd97}:		p = 14'd4559;
            {7'd47,7'd98}:		p = 14'd4606;
            {7'd47,7'd99}:		p = 14'd4653;
            {7'd47,7'd100}:		p = 14'd4700;
            {7'd47,7'd101}:		p = 14'd4747;
            {7'd47,7'd102}:		p = 14'd4794;
            {7'd47,7'd103}:		p = 14'd4841;
            {7'd47,7'd104}:		p = 14'd4888;
            {7'd47,7'd105}:		p = 14'd4935;
            {7'd47,7'd106}:		p = 14'd4982;
            {7'd47,7'd107}:		p = 14'd5029;
            {7'd47,7'd108}:		p = 14'd5076;
            {7'd47,7'd109}:		p = 14'd5123;
            {7'd47,7'd110}:		p = 14'd5170;
            {7'd47,7'd111}:		p = 14'd5217;
            {7'd47,7'd112}:		p = 14'd5264;
            {7'd47,7'd113}:		p = 14'd5311;
            {7'd47,7'd114}:		p = 14'd5358;
            {7'd47,7'd115}:		p = 14'd5405;
            {7'd47,7'd116}:		p = 14'd5452;
            {7'd47,7'd117}:		p = 14'd5499;
            {7'd47,7'd118}:		p = 14'd5546;
            {7'd47,7'd119}:		p = 14'd5593;
            {7'd47,7'd120}:		p = 14'd5640;
            {7'd47,7'd121}:		p = 14'd5687;
            {7'd47,7'd122}:		p = 14'd5734;
            {7'd47,7'd123}:		p = 14'd5781;
            {7'd47,7'd124}:		p = 14'd5828;
            {7'd47,7'd125}:		p = 14'd5875;
            {7'd47,7'd126}:		p = 14'd5922;
            {7'd47,7'd127}:		p = 14'd5969;
            {7'd48,7'd0}:		p = 14'd0;
            {7'd48,7'd1}:		p = 14'd48;
            {7'd48,7'd2}:		p = 14'd96;
            {7'd48,7'd3}:		p = 14'd144;
            {7'd48,7'd4}:		p = 14'd192;
            {7'd48,7'd5}:		p = 14'd240;
            {7'd48,7'd6}:		p = 14'd288;
            {7'd48,7'd7}:		p = 14'd336;
            {7'd48,7'd8}:		p = 14'd384;
            {7'd48,7'd9}:		p = 14'd432;
            {7'd48,7'd10}:		p = 14'd480;
            {7'd48,7'd11}:		p = 14'd528;
            {7'd48,7'd12}:		p = 14'd576;
            {7'd48,7'd13}:		p = 14'd624;
            {7'd48,7'd14}:		p = 14'd672;
            {7'd48,7'd15}:		p = 14'd720;
            {7'd48,7'd16}:		p = 14'd768;
            {7'd48,7'd17}:		p = 14'd816;
            {7'd48,7'd18}:		p = 14'd864;
            {7'd48,7'd19}:		p = 14'd912;
            {7'd48,7'd20}:		p = 14'd960;
            {7'd48,7'd21}:		p = 14'd1008;
            {7'd48,7'd22}:		p = 14'd1056;
            {7'd48,7'd23}:		p = 14'd1104;
            {7'd48,7'd24}:		p = 14'd1152;
            {7'd48,7'd25}:		p = 14'd1200;
            {7'd48,7'd26}:		p = 14'd1248;
            {7'd48,7'd27}:		p = 14'd1296;
            {7'd48,7'd28}:		p = 14'd1344;
            {7'd48,7'd29}:		p = 14'd1392;
            {7'd48,7'd30}:		p = 14'd1440;
            {7'd48,7'd31}:		p = 14'd1488;
            {7'd48,7'd32}:		p = 14'd1536;
            {7'd48,7'd33}:		p = 14'd1584;
            {7'd48,7'd34}:		p = 14'd1632;
            {7'd48,7'd35}:		p = 14'd1680;
            {7'd48,7'd36}:		p = 14'd1728;
            {7'd48,7'd37}:		p = 14'd1776;
            {7'd48,7'd38}:		p = 14'd1824;
            {7'd48,7'd39}:		p = 14'd1872;
            {7'd48,7'd40}:		p = 14'd1920;
            {7'd48,7'd41}:		p = 14'd1968;
            {7'd48,7'd42}:		p = 14'd2016;
            {7'd48,7'd43}:		p = 14'd2064;
            {7'd48,7'd44}:		p = 14'd2112;
            {7'd48,7'd45}:		p = 14'd2160;
            {7'd48,7'd46}:		p = 14'd2208;
            {7'd48,7'd47}:		p = 14'd2256;
            {7'd48,7'd48}:		p = 14'd2304;
            {7'd48,7'd49}:		p = 14'd2352;
            {7'd48,7'd50}:		p = 14'd2400;
            {7'd48,7'd51}:		p = 14'd2448;
            {7'd48,7'd52}:		p = 14'd2496;
            {7'd48,7'd53}:		p = 14'd2544;
            {7'd48,7'd54}:		p = 14'd2592;
            {7'd48,7'd55}:		p = 14'd2640;
            {7'd48,7'd56}:		p = 14'd2688;
            {7'd48,7'd57}:		p = 14'd2736;
            {7'd48,7'd58}:		p = 14'd2784;
            {7'd48,7'd59}:		p = 14'd2832;
            {7'd48,7'd60}:		p = 14'd2880;
            {7'd48,7'd61}:		p = 14'd2928;
            {7'd48,7'd62}:		p = 14'd2976;
            {7'd48,7'd63}:		p = 14'd3024;
            {7'd48,7'd64}:		p = 14'd3072;
            {7'd48,7'd65}:		p = 14'd3120;
            {7'd48,7'd66}:		p = 14'd3168;
            {7'd48,7'd67}:		p = 14'd3216;
            {7'd48,7'd68}:		p = 14'd3264;
            {7'd48,7'd69}:		p = 14'd3312;
            {7'd48,7'd70}:		p = 14'd3360;
            {7'd48,7'd71}:		p = 14'd3408;
            {7'd48,7'd72}:		p = 14'd3456;
            {7'd48,7'd73}:		p = 14'd3504;
            {7'd48,7'd74}:		p = 14'd3552;
            {7'd48,7'd75}:		p = 14'd3600;
            {7'd48,7'd76}:		p = 14'd3648;
            {7'd48,7'd77}:		p = 14'd3696;
            {7'd48,7'd78}:		p = 14'd3744;
            {7'd48,7'd79}:		p = 14'd3792;
            {7'd48,7'd80}:		p = 14'd3840;
            {7'd48,7'd81}:		p = 14'd3888;
            {7'd48,7'd82}:		p = 14'd3936;
            {7'd48,7'd83}:		p = 14'd3984;
            {7'd48,7'd84}:		p = 14'd4032;
            {7'd48,7'd85}:		p = 14'd4080;
            {7'd48,7'd86}:		p = 14'd4128;
            {7'd48,7'd87}:		p = 14'd4176;
            {7'd48,7'd88}:		p = 14'd4224;
            {7'd48,7'd89}:		p = 14'd4272;
            {7'd48,7'd90}:		p = 14'd4320;
            {7'd48,7'd91}:		p = 14'd4368;
            {7'd48,7'd92}:		p = 14'd4416;
            {7'd48,7'd93}:		p = 14'd4464;
            {7'd48,7'd94}:		p = 14'd4512;
            {7'd48,7'd95}:		p = 14'd4560;
            {7'd48,7'd96}:		p = 14'd4608;
            {7'd48,7'd97}:		p = 14'd4656;
            {7'd48,7'd98}:		p = 14'd4704;
            {7'd48,7'd99}:		p = 14'd4752;
            {7'd48,7'd100}:		p = 14'd4800;
            {7'd48,7'd101}:		p = 14'd4848;
            {7'd48,7'd102}:		p = 14'd4896;
            {7'd48,7'd103}:		p = 14'd4944;
            {7'd48,7'd104}:		p = 14'd4992;
            {7'd48,7'd105}:		p = 14'd5040;
            {7'd48,7'd106}:		p = 14'd5088;
            {7'd48,7'd107}:		p = 14'd5136;
            {7'd48,7'd108}:		p = 14'd5184;
            {7'd48,7'd109}:		p = 14'd5232;
            {7'd48,7'd110}:		p = 14'd5280;
            {7'd48,7'd111}:		p = 14'd5328;
            {7'd48,7'd112}:		p = 14'd5376;
            {7'd48,7'd113}:		p = 14'd5424;
            {7'd48,7'd114}:		p = 14'd5472;
            {7'd48,7'd115}:		p = 14'd5520;
            {7'd48,7'd116}:		p = 14'd5568;
            {7'd48,7'd117}:		p = 14'd5616;
            {7'd48,7'd118}:		p = 14'd5664;
            {7'd48,7'd119}:		p = 14'd5712;
            {7'd48,7'd120}:		p = 14'd5760;
            {7'd48,7'd121}:		p = 14'd5808;
            {7'd48,7'd122}:		p = 14'd5856;
            {7'd48,7'd123}:		p = 14'd5904;
            {7'd48,7'd124}:		p = 14'd5952;
            {7'd48,7'd125}:		p = 14'd6000;
            {7'd48,7'd126}:		p = 14'd6048;
            {7'd48,7'd127}:		p = 14'd6096;
            {7'd49,7'd0}:		p = 14'd0;
            {7'd49,7'd1}:		p = 14'd49;
            {7'd49,7'd2}:		p = 14'd98;
            {7'd49,7'd3}:		p = 14'd147;
            {7'd49,7'd4}:		p = 14'd196;
            {7'd49,7'd5}:		p = 14'd245;
            {7'd49,7'd6}:		p = 14'd294;
            {7'd49,7'd7}:		p = 14'd343;
            {7'd49,7'd8}:		p = 14'd392;
            {7'd49,7'd9}:		p = 14'd441;
            {7'd49,7'd10}:		p = 14'd490;
            {7'd49,7'd11}:		p = 14'd539;
            {7'd49,7'd12}:		p = 14'd588;
            {7'd49,7'd13}:		p = 14'd637;
            {7'd49,7'd14}:		p = 14'd686;
            {7'd49,7'd15}:		p = 14'd735;
            {7'd49,7'd16}:		p = 14'd784;
            {7'd49,7'd17}:		p = 14'd833;
            {7'd49,7'd18}:		p = 14'd882;
            {7'd49,7'd19}:		p = 14'd931;
            {7'd49,7'd20}:		p = 14'd980;
            {7'd49,7'd21}:		p = 14'd1029;
            {7'd49,7'd22}:		p = 14'd1078;
            {7'd49,7'd23}:		p = 14'd1127;
            {7'd49,7'd24}:		p = 14'd1176;
            {7'd49,7'd25}:		p = 14'd1225;
            {7'd49,7'd26}:		p = 14'd1274;
            {7'd49,7'd27}:		p = 14'd1323;
            {7'd49,7'd28}:		p = 14'd1372;
            {7'd49,7'd29}:		p = 14'd1421;
            {7'd49,7'd30}:		p = 14'd1470;
            {7'd49,7'd31}:		p = 14'd1519;
            {7'd49,7'd32}:		p = 14'd1568;
            {7'd49,7'd33}:		p = 14'd1617;
            {7'd49,7'd34}:		p = 14'd1666;
            {7'd49,7'd35}:		p = 14'd1715;
            {7'd49,7'd36}:		p = 14'd1764;
            {7'd49,7'd37}:		p = 14'd1813;
            {7'd49,7'd38}:		p = 14'd1862;
            {7'd49,7'd39}:		p = 14'd1911;
            {7'd49,7'd40}:		p = 14'd1960;
            {7'd49,7'd41}:		p = 14'd2009;
            {7'd49,7'd42}:		p = 14'd2058;
            {7'd49,7'd43}:		p = 14'd2107;
            {7'd49,7'd44}:		p = 14'd2156;
            {7'd49,7'd45}:		p = 14'd2205;
            {7'd49,7'd46}:		p = 14'd2254;
            {7'd49,7'd47}:		p = 14'd2303;
            {7'd49,7'd48}:		p = 14'd2352;
            {7'd49,7'd49}:		p = 14'd2401;
            {7'd49,7'd50}:		p = 14'd2450;
            {7'd49,7'd51}:		p = 14'd2499;
            {7'd49,7'd52}:		p = 14'd2548;
            {7'd49,7'd53}:		p = 14'd2597;
            {7'd49,7'd54}:		p = 14'd2646;
            {7'd49,7'd55}:		p = 14'd2695;
            {7'd49,7'd56}:		p = 14'd2744;
            {7'd49,7'd57}:		p = 14'd2793;
            {7'd49,7'd58}:		p = 14'd2842;
            {7'd49,7'd59}:		p = 14'd2891;
            {7'd49,7'd60}:		p = 14'd2940;
            {7'd49,7'd61}:		p = 14'd2989;
            {7'd49,7'd62}:		p = 14'd3038;
            {7'd49,7'd63}:		p = 14'd3087;
            {7'd49,7'd64}:		p = 14'd3136;
            {7'd49,7'd65}:		p = 14'd3185;
            {7'd49,7'd66}:		p = 14'd3234;
            {7'd49,7'd67}:		p = 14'd3283;
            {7'd49,7'd68}:		p = 14'd3332;
            {7'd49,7'd69}:		p = 14'd3381;
            {7'd49,7'd70}:		p = 14'd3430;
            {7'd49,7'd71}:		p = 14'd3479;
            {7'd49,7'd72}:		p = 14'd3528;
            {7'd49,7'd73}:		p = 14'd3577;
            {7'd49,7'd74}:		p = 14'd3626;
            {7'd49,7'd75}:		p = 14'd3675;
            {7'd49,7'd76}:		p = 14'd3724;
            {7'd49,7'd77}:		p = 14'd3773;
            {7'd49,7'd78}:		p = 14'd3822;
            {7'd49,7'd79}:		p = 14'd3871;
            {7'd49,7'd80}:		p = 14'd3920;
            {7'd49,7'd81}:		p = 14'd3969;
            {7'd49,7'd82}:		p = 14'd4018;
            {7'd49,7'd83}:		p = 14'd4067;
            {7'd49,7'd84}:		p = 14'd4116;
            {7'd49,7'd85}:		p = 14'd4165;
            {7'd49,7'd86}:		p = 14'd4214;
            {7'd49,7'd87}:		p = 14'd4263;
            {7'd49,7'd88}:		p = 14'd4312;
            {7'd49,7'd89}:		p = 14'd4361;
            {7'd49,7'd90}:		p = 14'd4410;
            {7'd49,7'd91}:		p = 14'd4459;
            {7'd49,7'd92}:		p = 14'd4508;
            {7'd49,7'd93}:		p = 14'd4557;
            {7'd49,7'd94}:		p = 14'd4606;
            {7'd49,7'd95}:		p = 14'd4655;
            {7'd49,7'd96}:		p = 14'd4704;
            {7'd49,7'd97}:		p = 14'd4753;
            {7'd49,7'd98}:		p = 14'd4802;
            {7'd49,7'd99}:		p = 14'd4851;
            {7'd49,7'd100}:		p = 14'd4900;
            {7'd49,7'd101}:		p = 14'd4949;
            {7'd49,7'd102}:		p = 14'd4998;
            {7'd49,7'd103}:		p = 14'd5047;
            {7'd49,7'd104}:		p = 14'd5096;
            {7'd49,7'd105}:		p = 14'd5145;
            {7'd49,7'd106}:		p = 14'd5194;
            {7'd49,7'd107}:		p = 14'd5243;
            {7'd49,7'd108}:		p = 14'd5292;
            {7'd49,7'd109}:		p = 14'd5341;
            {7'd49,7'd110}:		p = 14'd5390;
            {7'd49,7'd111}:		p = 14'd5439;
            {7'd49,7'd112}:		p = 14'd5488;
            {7'd49,7'd113}:		p = 14'd5537;
            {7'd49,7'd114}:		p = 14'd5586;
            {7'd49,7'd115}:		p = 14'd5635;
            {7'd49,7'd116}:		p = 14'd5684;
            {7'd49,7'd117}:		p = 14'd5733;
            {7'd49,7'd118}:		p = 14'd5782;
            {7'd49,7'd119}:		p = 14'd5831;
            {7'd49,7'd120}:		p = 14'd5880;
            {7'd49,7'd121}:		p = 14'd5929;
            {7'd49,7'd122}:		p = 14'd5978;
            {7'd49,7'd123}:		p = 14'd6027;
            {7'd49,7'd124}:		p = 14'd6076;
            {7'd49,7'd125}:		p = 14'd6125;
            {7'd49,7'd126}:		p = 14'd6174;
            {7'd49,7'd127}:		p = 14'd6223;
            {7'd50,7'd0}:		p = 14'd0;
            {7'd50,7'd1}:		p = 14'd50;
            {7'd50,7'd2}:		p = 14'd100;
            {7'd50,7'd3}:		p = 14'd150;
            {7'd50,7'd4}:		p = 14'd200;
            {7'd50,7'd5}:		p = 14'd250;
            {7'd50,7'd6}:		p = 14'd300;
            {7'd50,7'd7}:		p = 14'd350;
            {7'd50,7'd8}:		p = 14'd400;
            {7'd50,7'd9}:		p = 14'd450;
            {7'd50,7'd10}:		p = 14'd500;
            {7'd50,7'd11}:		p = 14'd550;
            {7'd50,7'd12}:		p = 14'd600;
            {7'd50,7'd13}:		p = 14'd650;
            {7'd50,7'd14}:		p = 14'd700;
            {7'd50,7'd15}:		p = 14'd750;
            {7'd50,7'd16}:		p = 14'd800;
            {7'd50,7'd17}:		p = 14'd850;
            {7'd50,7'd18}:		p = 14'd900;
            {7'd50,7'd19}:		p = 14'd950;
            {7'd50,7'd20}:		p = 14'd1000;
            {7'd50,7'd21}:		p = 14'd1050;
            {7'd50,7'd22}:		p = 14'd1100;
            {7'd50,7'd23}:		p = 14'd1150;
            {7'd50,7'd24}:		p = 14'd1200;
            {7'd50,7'd25}:		p = 14'd1250;
            {7'd50,7'd26}:		p = 14'd1300;
            {7'd50,7'd27}:		p = 14'd1350;
            {7'd50,7'd28}:		p = 14'd1400;
            {7'd50,7'd29}:		p = 14'd1450;
            {7'd50,7'd30}:		p = 14'd1500;
            {7'd50,7'd31}:		p = 14'd1550;
            {7'd50,7'd32}:		p = 14'd1600;
            {7'd50,7'd33}:		p = 14'd1650;
            {7'd50,7'd34}:		p = 14'd1700;
            {7'd50,7'd35}:		p = 14'd1750;
            {7'd50,7'd36}:		p = 14'd1800;
            {7'd50,7'd37}:		p = 14'd1850;
            {7'd50,7'd38}:		p = 14'd1900;
            {7'd50,7'd39}:		p = 14'd1950;
            {7'd50,7'd40}:		p = 14'd2000;
            {7'd50,7'd41}:		p = 14'd2050;
            {7'd50,7'd42}:		p = 14'd2100;
            {7'd50,7'd43}:		p = 14'd2150;
            {7'd50,7'd44}:		p = 14'd2200;
            {7'd50,7'd45}:		p = 14'd2250;
            {7'd50,7'd46}:		p = 14'd2300;
            {7'd50,7'd47}:		p = 14'd2350;
            {7'd50,7'd48}:		p = 14'd2400;
            {7'd50,7'd49}:		p = 14'd2450;
            {7'd50,7'd50}:		p = 14'd2500;
            {7'd50,7'd51}:		p = 14'd2550;
            {7'd50,7'd52}:		p = 14'd2600;
            {7'd50,7'd53}:		p = 14'd2650;
            {7'd50,7'd54}:		p = 14'd2700;
            {7'd50,7'd55}:		p = 14'd2750;
            {7'd50,7'd56}:		p = 14'd2800;
            {7'd50,7'd57}:		p = 14'd2850;
            {7'd50,7'd58}:		p = 14'd2900;
            {7'd50,7'd59}:		p = 14'd2950;
            {7'd50,7'd60}:		p = 14'd3000;
            {7'd50,7'd61}:		p = 14'd3050;
            {7'd50,7'd62}:		p = 14'd3100;
            {7'd50,7'd63}:		p = 14'd3150;
            {7'd50,7'd64}:		p = 14'd3200;
            {7'd50,7'd65}:		p = 14'd3250;
            {7'd50,7'd66}:		p = 14'd3300;
            {7'd50,7'd67}:		p = 14'd3350;
            {7'd50,7'd68}:		p = 14'd3400;
            {7'd50,7'd69}:		p = 14'd3450;
            {7'd50,7'd70}:		p = 14'd3500;
            {7'd50,7'd71}:		p = 14'd3550;
            {7'd50,7'd72}:		p = 14'd3600;
            {7'd50,7'd73}:		p = 14'd3650;
            {7'd50,7'd74}:		p = 14'd3700;
            {7'd50,7'd75}:		p = 14'd3750;
            {7'd50,7'd76}:		p = 14'd3800;
            {7'd50,7'd77}:		p = 14'd3850;
            {7'd50,7'd78}:		p = 14'd3900;
            {7'd50,7'd79}:		p = 14'd3950;
            {7'd50,7'd80}:		p = 14'd4000;
            {7'd50,7'd81}:		p = 14'd4050;
            {7'd50,7'd82}:		p = 14'd4100;
            {7'd50,7'd83}:		p = 14'd4150;
            {7'd50,7'd84}:		p = 14'd4200;
            {7'd50,7'd85}:		p = 14'd4250;
            {7'd50,7'd86}:		p = 14'd4300;
            {7'd50,7'd87}:		p = 14'd4350;
            {7'd50,7'd88}:		p = 14'd4400;
            {7'd50,7'd89}:		p = 14'd4450;
            {7'd50,7'd90}:		p = 14'd4500;
            {7'd50,7'd91}:		p = 14'd4550;
            {7'd50,7'd92}:		p = 14'd4600;
            {7'd50,7'd93}:		p = 14'd4650;
            {7'd50,7'd94}:		p = 14'd4700;
            {7'd50,7'd95}:		p = 14'd4750;
            {7'd50,7'd96}:		p = 14'd4800;
            {7'd50,7'd97}:		p = 14'd4850;
            {7'd50,7'd98}:		p = 14'd4900;
            {7'd50,7'd99}:		p = 14'd4950;
            {7'd50,7'd100}:		p = 14'd5000;
            {7'd50,7'd101}:		p = 14'd5050;
            {7'd50,7'd102}:		p = 14'd5100;
            {7'd50,7'd103}:		p = 14'd5150;
            {7'd50,7'd104}:		p = 14'd5200;
            {7'd50,7'd105}:		p = 14'd5250;
            {7'd50,7'd106}:		p = 14'd5300;
            {7'd50,7'd107}:		p = 14'd5350;
            {7'd50,7'd108}:		p = 14'd5400;
            {7'd50,7'd109}:		p = 14'd5450;
            {7'd50,7'd110}:		p = 14'd5500;
            {7'd50,7'd111}:		p = 14'd5550;
            {7'd50,7'd112}:		p = 14'd5600;
            {7'd50,7'd113}:		p = 14'd5650;
            {7'd50,7'd114}:		p = 14'd5700;
            {7'd50,7'd115}:		p = 14'd5750;
            {7'd50,7'd116}:		p = 14'd5800;
            {7'd50,7'd117}:		p = 14'd5850;
            {7'd50,7'd118}:		p = 14'd5900;
            {7'd50,7'd119}:		p = 14'd5950;
            {7'd50,7'd120}:		p = 14'd6000;
            {7'd50,7'd121}:		p = 14'd6050;
            {7'd50,7'd122}:		p = 14'd6100;
            {7'd50,7'd123}:		p = 14'd6150;
            {7'd50,7'd124}:		p = 14'd6200;
            {7'd50,7'd125}:		p = 14'd6250;
            {7'd50,7'd126}:		p = 14'd6300;
            {7'd50,7'd127}:		p = 14'd6350;
            {7'd51,7'd0}:		p = 14'd0;
            {7'd51,7'd1}:		p = 14'd51;
            {7'd51,7'd2}:		p = 14'd102;
            {7'd51,7'd3}:		p = 14'd153;
            {7'd51,7'd4}:		p = 14'd204;
            {7'd51,7'd5}:		p = 14'd255;
            {7'd51,7'd6}:		p = 14'd306;
            {7'd51,7'd7}:		p = 14'd357;
            {7'd51,7'd8}:		p = 14'd408;
            {7'd51,7'd9}:		p = 14'd459;
            {7'd51,7'd10}:		p = 14'd510;
            {7'd51,7'd11}:		p = 14'd561;
            {7'd51,7'd12}:		p = 14'd612;
            {7'd51,7'd13}:		p = 14'd663;
            {7'd51,7'd14}:		p = 14'd714;
            {7'd51,7'd15}:		p = 14'd765;
            {7'd51,7'd16}:		p = 14'd816;
            {7'd51,7'd17}:		p = 14'd867;
            {7'd51,7'd18}:		p = 14'd918;
            {7'd51,7'd19}:		p = 14'd969;
            {7'd51,7'd20}:		p = 14'd1020;
            {7'd51,7'd21}:		p = 14'd1071;
            {7'd51,7'd22}:		p = 14'd1122;
            {7'd51,7'd23}:		p = 14'd1173;
            {7'd51,7'd24}:		p = 14'd1224;
            {7'd51,7'd25}:		p = 14'd1275;
            {7'd51,7'd26}:		p = 14'd1326;
            {7'd51,7'd27}:		p = 14'd1377;
            {7'd51,7'd28}:		p = 14'd1428;
            {7'd51,7'd29}:		p = 14'd1479;
            {7'd51,7'd30}:		p = 14'd1530;
            {7'd51,7'd31}:		p = 14'd1581;
            {7'd51,7'd32}:		p = 14'd1632;
            {7'd51,7'd33}:		p = 14'd1683;
            {7'd51,7'd34}:		p = 14'd1734;
            {7'd51,7'd35}:		p = 14'd1785;
            {7'd51,7'd36}:		p = 14'd1836;
            {7'd51,7'd37}:		p = 14'd1887;
            {7'd51,7'd38}:		p = 14'd1938;
            {7'd51,7'd39}:		p = 14'd1989;
            {7'd51,7'd40}:		p = 14'd2040;
            {7'd51,7'd41}:		p = 14'd2091;
            {7'd51,7'd42}:		p = 14'd2142;
            {7'd51,7'd43}:		p = 14'd2193;
            {7'd51,7'd44}:		p = 14'd2244;
            {7'd51,7'd45}:		p = 14'd2295;
            {7'd51,7'd46}:		p = 14'd2346;
            {7'd51,7'd47}:		p = 14'd2397;
            {7'd51,7'd48}:		p = 14'd2448;
            {7'd51,7'd49}:		p = 14'd2499;
            {7'd51,7'd50}:		p = 14'd2550;
            {7'd51,7'd51}:		p = 14'd2601;
            {7'd51,7'd52}:		p = 14'd2652;
            {7'd51,7'd53}:		p = 14'd2703;
            {7'd51,7'd54}:		p = 14'd2754;
            {7'd51,7'd55}:		p = 14'd2805;
            {7'd51,7'd56}:		p = 14'd2856;
            {7'd51,7'd57}:		p = 14'd2907;
            {7'd51,7'd58}:		p = 14'd2958;
            {7'd51,7'd59}:		p = 14'd3009;
            {7'd51,7'd60}:		p = 14'd3060;
            {7'd51,7'd61}:		p = 14'd3111;
            {7'd51,7'd62}:		p = 14'd3162;
            {7'd51,7'd63}:		p = 14'd3213;
            {7'd51,7'd64}:		p = 14'd3264;
            {7'd51,7'd65}:		p = 14'd3315;
            {7'd51,7'd66}:		p = 14'd3366;
            {7'd51,7'd67}:		p = 14'd3417;
            {7'd51,7'd68}:		p = 14'd3468;
            {7'd51,7'd69}:		p = 14'd3519;
            {7'd51,7'd70}:		p = 14'd3570;
            {7'd51,7'd71}:		p = 14'd3621;
            {7'd51,7'd72}:		p = 14'd3672;
            {7'd51,7'd73}:		p = 14'd3723;
            {7'd51,7'd74}:		p = 14'd3774;
            {7'd51,7'd75}:		p = 14'd3825;
            {7'd51,7'd76}:		p = 14'd3876;
            {7'd51,7'd77}:		p = 14'd3927;
            {7'd51,7'd78}:		p = 14'd3978;
            {7'd51,7'd79}:		p = 14'd4029;
            {7'd51,7'd80}:		p = 14'd4080;
            {7'd51,7'd81}:		p = 14'd4131;
            {7'd51,7'd82}:		p = 14'd4182;
            {7'd51,7'd83}:		p = 14'd4233;
            {7'd51,7'd84}:		p = 14'd4284;
            {7'd51,7'd85}:		p = 14'd4335;
            {7'd51,7'd86}:		p = 14'd4386;
            {7'd51,7'd87}:		p = 14'd4437;
            {7'd51,7'd88}:		p = 14'd4488;
            {7'd51,7'd89}:		p = 14'd4539;
            {7'd51,7'd90}:		p = 14'd4590;
            {7'd51,7'd91}:		p = 14'd4641;
            {7'd51,7'd92}:		p = 14'd4692;
            {7'd51,7'd93}:		p = 14'd4743;
            {7'd51,7'd94}:		p = 14'd4794;
            {7'd51,7'd95}:		p = 14'd4845;
            {7'd51,7'd96}:		p = 14'd4896;
            {7'd51,7'd97}:		p = 14'd4947;
            {7'd51,7'd98}:		p = 14'd4998;
            {7'd51,7'd99}:		p = 14'd5049;
            {7'd51,7'd100}:		p = 14'd5100;
            {7'd51,7'd101}:		p = 14'd5151;
            {7'd51,7'd102}:		p = 14'd5202;
            {7'd51,7'd103}:		p = 14'd5253;
            {7'd51,7'd104}:		p = 14'd5304;
            {7'd51,7'd105}:		p = 14'd5355;
            {7'd51,7'd106}:		p = 14'd5406;
            {7'd51,7'd107}:		p = 14'd5457;
            {7'd51,7'd108}:		p = 14'd5508;
            {7'd51,7'd109}:		p = 14'd5559;
            {7'd51,7'd110}:		p = 14'd5610;
            {7'd51,7'd111}:		p = 14'd5661;
            {7'd51,7'd112}:		p = 14'd5712;
            {7'd51,7'd113}:		p = 14'd5763;
            {7'd51,7'd114}:		p = 14'd5814;
            {7'd51,7'd115}:		p = 14'd5865;
            {7'd51,7'd116}:		p = 14'd5916;
            {7'd51,7'd117}:		p = 14'd5967;
            {7'd51,7'd118}:		p = 14'd6018;
            {7'd51,7'd119}:		p = 14'd6069;
            {7'd51,7'd120}:		p = 14'd6120;
            {7'd51,7'd121}:		p = 14'd6171;
            {7'd51,7'd122}:		p = 14'd6222;
            {7'd51,7'd123}:		p = 14'd6273;
            {7'd51,7'd124}:		p = 14'd6324;
            {7'd51,7'd125}:		p = 14'd6375;
            {7'd51,7'd126}:		p = 14'd6426;
            {7'd51,7'd127}:		p = 14'd6477;
            {7'd52,7'd0}:		p = 14'd0;
            {7'd52,7'd1}:		p = 14'd52;
            {7'd52,7'd2}:		p = 14'd104;
            {7'd52,7'd3}:		p = 14'd156;
            {7'd52,7'd4}:		p = 14'd208;
            {7'd52,7'd5}:		p = 14'd260;
            {7'd52,7'd6}:		p = 14'd312;
            {7'd52,7'd7}:		p = 14'd364;
            {7'd52,7'd8}:		p = 14'd416;
            {7'd52,7'd9}:		p = 14'd468;
            {7'd52,7'd10}:		p = 14'd520;
            {7'd52,7'd11}:		p = 14'd572;
            {7'd52,7'd12}:		p = 14'd624;
            {7'd52,7'd13}:		p = 14'd676;
            {7'd52,7'd14}:		p = 14'd728;
            {7'd52,7'd15}:		p = 14'd780;
            {7'd52,7'd16}:		p = 14'd832;
            {7'd52,7'd17}:		p = 14'd884;
            {7'd52,7'd18}:		p = 14'd936;
            {7'd52,7'd19}:		p = 14'd988;
            {7'd52,7'd20}:		p = 14'd1040;
            {7'd52,7'd21}:		p = 14'd1092;
            {7'd52,7'd22}:		p = 14'd1144;
            {7'd52,7'd23}:		p = 14'd1196;
            {7'd52,7'd24}:		p = 14'd1248;
            {7'd52,7'd25}:		p = 14'd1300;
            {7'd52,7'd26}:		p = 14'd1352;
            {7'd52,7'd27}:		p = 14'd1404;
            {7'd52,7'd28}:		p = 14'd1456;
            {7'd52,7'd29}:		p = 14'd1508;
            {7'd52,7'd30}:		p = 14'd1560;
            {7'd52,7'd31}:		p = 14'd1612;
            {7'd52,7'd32}:		p = 14'd1664;
            {7'd52,7'd33}:		p = 14'd1716;
            {7'd52,7'd34}:		p = 14'd1768;
            {7'd52,7'd35}:		p = 14'd1820;
            {7'd52,7'd36}:		p = 14'd1872;
            {7'd52,7'd37}:		p = 14'd1924;
            {7'd52,7'd38}:		p = 14'd1976;
            {7'd52,7'd39}:		p = 14'd2028;
            {7'd52,7'd40}:		p = 14'd2080;
            {7'd52,7'd41}:		p = 14'd2132;
            {7'd52,7'd42}:		p = 14'd2184;
            {7'd52,7'd43}:		p = 14'd2236;
            {7'd52,7'd44}:		p = 14'd2288;
            {7'd52,7'd45}:		p = 14'd2340;
            {7'd52,7'd46}:		p = 14'd2392;
            {7'd52,7'd47}:		p = 14'd2444;
            {7'd52,7'd48}:		p = 14'd2496;
            {7'd52,7'd49}:		p = 14'd2548;
            {7'd52,7'd50}:		p = 14'd2600;
            {7'd52,7'd51}:		p = 14'd2652;
            {7'd52,7'd52}:		p = 14'd2704;
            {7'd52,7'd53}:		p = 14'd2756;
            {7'd52,7'd54}:		p = 14'd2808;
            {7'd52,7'd55}:		p = 14'd2860;
            {7'd52,7'd56}:		p = 14'd2912;
            {7'd52,7'd57}:		p = 14'd2964;
            {7'd52,7'd58}:		p = 14'd3016;
            {7'd52,7'd59}:		p = 14'd3068;
            {7'd52,7'd60}:		p = 14'd3120;
            {7'd52,7'd61}:		p = 14'd3172;
            {7'd52,7'd62}:		p = 14'd3224;
            {7'd52,7'd63}:		p = 14'd3276;
            {7'd52,7'd64}:		p = 14'd3328;
            {7'd52,7'd65}:		p = 14'd3380;
            {7'd52,7'd66}:		p = 14'd3432;
            {7'd52,7'd67}:		p = 14'd3484;
            {7'd52,7'd68}:		p = 14'd3536;
            {7'd52,7'd69}:		p = 14'd3588;
            {7'd52,7'd70}:		p = 14'd3640;
            {7'd52,7'd71}:		p = 14'd3692;
            {7'd52,7'd72}:		p = 14'd3744;
            {7'd52,7'd73}:		p = 14'd3796;
            {7'd52,7'd74}:		p = 14'd3848;
            {7'd52,7'd75}:		p = 14'd3900;
            {7'd52,7'd76}:		p = 14'd3952;
            {7'd52,7'd77}:		p = 14'd4004;
            {7'd52,7'd78}:		p = 14'd4056;
            {7'd52,7'd79}:		p = 14'd4108;
            {7'd52,7'd80}:		p = 14'd4160;
            {7'd52,7'd81}:		p = 14'd4212;
            {7'd52,7'd82}:		p = 14'd4264;
            {7'd52,7'd83}:		p = 14'd4316;
            {7'd52,7'd84}:		p = 14'd4368;
            {7'd52,7'd85}:		p = 14'd4420;
            {7'd52,7'd86}:		p = 14'd4472;
            {7'd52,7'd87}:		p = 14'd4524;
            {7'd52,7'd88}:		p = 14'd4576;
            {7'd52,7'd89}:		p = 14'd4628;
            {7'd52,7'd90}:		p = 14'd4680;
            {7'd52,7'd91}:		p = 14'd4732;
            {7'd52,7'd92}:		p = 14'd4784;
            {7'd52,7'd93}:		p = 14'd4836;
            {7'd52,7'd94}:		p = 14'd4888;
            {7'd52,7'd95}:		p = 14'd4940;
            {7'd52,7'd96}:		p = 14'd4992;
            {7'd52,7'd97}:		p = 14'd5044;
            {7'd52,7'd98}:		p = 14'd5096;
            {7'd52,7'd99}:		p = 14'd5148;
            {7'd52,7'd100}:		p = 14'd5200;
            {7'd52,7'd101}:		p = 14'd5252;
            {7'd52,7'd102}:		p = 14'd5304;
            {7'd52,7'd103}:		p = 14'd5356;
            {7'd52,7'd104}:		p = 14'd5408;
            {7'd52,7'd105}:		p = 14'd5460;
            {7'd52,7'd106}:		p = 14'd5512;
            {7'd52,7'd107}:		p = 14'd5564;
            {7'd52,7'd108}:		p = 14'd5616;
            {7'd52,7'd109}:		p = 14'd5668;
            {7'd52,7'd110}:		p = 14'd5720;
            {7'd52,7'd111}:		p = 14'd5772;
            {7'd52,7'd112}:		p = 14'd5824;
            {7'd52,7'd113}:		p = 14'd5876;
            {7'd52,7'd114}:		p = 14'd5928;
            {7'd52,7'd115}:		p = 14'd5980;
            {7'd52,7'd116}:		p = 14'd6032;
            {7'd52,7'd117}:		p = 14'd6084;
            {7'd52,7'd118}:		p = 14'd6136;
            {7'd52,7'd119}:		p = 14'd6188;
            {7'd52,7'd120}:		p = 14'd6240;
            {7'd52,7'd121}:		p = 14'd6292;
            {7'd52,7'd122}:		p = 14'd6344;
            {7'd52,7'd123}:		p = 14'd6396;
            {7'd52,7'd124}:		p = 14'd6448;
            {7'd52,7'd125}:		p = 14'd6500;
            {7'd52,7'd126}:		p = 14'd6552;
            {7'd52,7'd127}:		p = 14'd6604;
            {7'd53,7'd0}:		p = 14'd0;
            {7'd53,7'd1}:		p = 14'd53;
            {7'd53,7'd2}:		p = 14'd106;
            {7'd53,7'd3}:		p = 14'd159;
            {7'd53,7'd4}:		p = 14'd212;
            {7'd53,7'd5}:		p = 14'd265;
            {7'd53,7'd6}:		p = 14'd318;
            {7'd53,7'd7}:		p = 14'd371;
            {7'd53,7'd8}:		p = 14'd424;
            {7'd53,7'd9}:		p = 14'd477;
            {7'd53,7'd10}:		p = 14'd530;
            {7'd53,7'd11}:		p = 14'd583;
            {7'd53,7'd12}:		p = 14'd636;
            {7'd53,7'd13}:		p = 14'd689;
            {7'd53,7'd14}:		p = 14'd742;
            {7'd53,7'd15}:		p = 14'd795;
            {7'd53,7'd16}:		p = 14'd848;
            {7'd53,7'd17}:		p = 14'd901;
            {7'd53,7'd18}:		p = 14'd954;
            {7'd53,7'd19}:		p = 14'd1007;
            {7'd53,7'd20}:		p = 14'd1060;
            {7'd53,7'd21}:		p = 14'd1113;
            {7'd53,7'd22}:		p = 14'd1166;
            {7'd53,7'd23}:		p = 14'd1219;
            {7'd53,7'd24}:		p = 14'd1272;
            {7'd53,7'd25}:		p = 14'd1325;
            {7'd53,7'd26}:		p = 14'd1378;
            {7'd53,7'd27}:		p = 14'd1431;
            {7'd53,7'd28}:		p = 14'd1484;
            {7'd53,7'd29}:		p = 14'd1537;
            {7'd53,7'd30}:		p = 14'd1590;
            {7'd53,7'd31}:		p = 14'd1643;
            {7'd53,7'd32}:		p = 14'd1696;
            {7'd53,7'd33}:		p = 14'd1749;
            {7'd53,7'd34}:		p = 14'd1802;
            {7'd53,7'd35}:		p = 14'd1855;
            {7'd53,7'd36}:		p = 14'd1908;
            {7'd53,7'd37}:		p = 14'd1961;
            {7'd53,7'd38}:		p = 14'd2014;
            {7'd53,7'd39}:		p = 14'd2067;
            {7'd53,7'd40}:		p = 14'd2120;
            {7'd53,7'd41}:		p = 14'd2173;
            {7'd53,7'd42}:		p = 14'd2226;
            {7'd53,7'd43}:		p = 14'd2279;
            {7'd53,7'd44}:		p = 14'd2332;
            {7'd53,7'd45}:		p = 14'd2385;
            {7'd53,7'd46}:		p = 14'd2438;
            {7'd53,7'd47}:		p = 14'd2491;
            {7'd53,7'd48}:		p = 14'd2544;
            {7'd53,7'd49}:		p = 14'd2597;
            {7'd53,7'd50}:		p = 14'd2650;
            {7'd53,7'd51}:		p = 14'd2703;
            {7'd53,7'd52}:		p = 14'd2756;
            {7'd53,7'd53}:		p = 14'd2809;
            {7'd53,7'd54}:		p = 14'd2862;
            {7'd53,7'd55}:		p = 14'd2915;
            {7'd53,7'd56}:		p = 14'd2968;
            {7'd53,7'd57}:		p = 14'd3021;
            {7'd53,7'd58}:		p = 14'd3074;
            {7'd53,7'd59}:		p = 14'd3127;
            {7'd53,7'd60}:		p = 14'd3180;
            {7'd53,7'd61}:		p = 14'd3233;
            {7'd53,7'd62}:		p = 14'd3286;
            {7'd53,7'd63}:		p = 14'd3339;
            {7'd53,7'd64}:		p = 14'd3392;
            {7'd53,7'd65}:		p = 14'd3445;
            {7'd53,7'd66}:		p = 14'd3498;
            {7'd53,7'd67}:		p = 14'd3551;
            {7'd53,7'd68}:		p = 14'd3604;
            {7'd53,7'd69}:		p = 14'd3657;
            {7'd53,7'd70}:		p = 14'd3710;
            {7'd53,7'd71}:		p = 14'd3763;
            {7'd53,7'd72}:		p = 14'd3816;
            {7'd53,7'd73}:		p = 14'd3869;
            {7'd53,7'd74}:		p = 14'd3922;
            {7'd53,7'd75}:		p = 14'd3975;
            {7'd53,7'd76}:		p = 14'd4028;
            {7'd53,7'd77}:		p = 14'd4081;
            {7'd53,7'd78}:		p = 14'd4134;
            {7'd53,7'd79}:		p = 14'd4187;
            {7'd53,7'd80}:		p = 14'd4240;
            {7'd53,7'd81}:		p = 14'd4293;
            {7'd53,7'd82}:		p = 14'd4346;
            {7'd53,7'd83}:		p = 14'd4399;
            {7'd53,7'd84}:		p = 14'd4452;
            {7'd53,7'd85}:		p = 14'd4505;
            {7'd53,7'd86}:		p = 14'd4558;
            {7'd53,7'd87}:		p = 14'd4611;
            {7'd53,7'd88}:		p = 14'd4664;
            {7'd53,7'd89}:		p = 14'd4717;
            {7'd53,7'd90}:		p = 14'd4770;
            {7'd53,7'd91}:		p = 14'd4823;
            {7'd53,7'd92}:		p = 14'd4876;
            {7'd53,7'd93}:		p = 14'd4929;
            {7'd53,7'd94}:		p = 14'd4982;
            {7'd53,7'd95}:		p = 14'd5035;
            {7'd53,7'd96}:		p = 14'd5088;
            {7'd53,7'd97}:		p = 14'd5141;
            {7'd53,7'd98}:		p = 14'd5194;
            {7'd53,7'd99}:		p = 14'd5247;
            {7'd53,7'd100}:		p = 14'd5300;
            {7'd53,7'd101}:		p = 14'd5353;
            {7'd53,7'd102}:		p = 14'd5406;
            {7'd53,7'd103}:		p = 14'd5459;
            {7'd53,7'd104}:		p = 14'd5512;
            {7'd53,7'd105}:		p = 14'd5565;
            {7'd53,7'd106}:		p = 14'd5618;
            {7'd53,7'd107}:		p = 14'd5671;
            {7'd53,7'd108}:		p = 14'd5724;
            {7'd53,7'd109}:		p = 14'd5777;
            {7'd53,7'd110}:		p = 14'd5830;
            {7'd53,7'd111}:		p = 14'd5883;
            {7'd53,7'd112}:		p = 14'd5936;
            {7'd53,7'd113}:		p = 14'd5989;
            {7'd53,7'd114}:		p = 14'd6042;
            {7'd53,7'd115}:		p = 14'd6095;
            {7'd53,7'd116}:		p = 14'd6148;
            {7'd53,7'd117}:		p = 14'd6201;
            {7'd53,7'd118}:		p = 14'd6254;
            {7'd53,7'd119}:		p = 14'd6307;
            {7'd53,7'd120}:		p = 14'd6360;
            {7'd53,7'd121}:		p = 14'd6413;
            {7'd53,7'd122}:		p = 14'd6466;
            {7'd53,7'd123}:		p = 14'd6519;
            {7'd53,7'd124}:		p = 14'd6572;
            {7'd53,7'd125}:		p = 14'd6625;
            {7'd53,7'd126}:		p = 14'd6678;
            {7'd53,7'd127}:		p = 14'd6731;
            {7'd54,7'd0}:		p = 14'd0;
            {7'd54,7'd1}:		p = 14'd54;
            {7'd54,7'd2}:		p = 14'd108;
            {7'd54,7'd3}:		p = 14'd162;
            {7'd54,7'd4}:		p = 14'd216;
            {7'd54,7'd5}:		p = 14'd270;
            {7'd54,7'd6}:		p = 14'd324;
            {7'd54,7'd7}:		p = 14'd378;
            {7'd54,7'd8}:		p = 14'd432;
            {7'd54,7'd9}:		p = 14'd486;
            {7'd54,7'd10}:		p = 14'd540;
            {7'd54,7'd11}:		p = 14'd594;
            {7'd54,7'd12}:		p = 14'd648;
            {7'd54,7'd13}:		p = 14'd702;
            {7'd54,7'd14}:		p = 14'd756;
            {7'd54,7'd15}:		p = 14'd810;
            {7'd54,7'd16}:		p = 14'd864;
            {7'd54,7'd17}:		p = 14'd918;
            {7'd54,7'd18}:		p = 14'd972;
            {7'd54,7'd19}:		p = 14'd1026;
            {7'd54,7'd20}:		p = 14'd1080;
            {7'd54,7'd21}:		p = 14'd1134;
            {7'd54,7'd22}:		p = 14'd1188;
            {7'd54,7'd23}:		p = 14'd1242;
            {7'd54,7'd24}:		p = 14'd1296;
            {7'd54,7'd25}:		p = 14'd1350;
            {7'd54,7'd26}:		p = 14'd1404;
            {7'd54,7'd27}:		p = 14'd1458;
            {7'd54,7'd28}:		p = 14'd1512;
            {7'd54,7'd29}:		p = 14'd1566;
            {7'd54,7'd30}:		p = 14'd1620;
            {7'd54,7'd31}:		p = 14'd1674;
            {7'd54,7'd32}:		p = 14'd1728;
            {7'd54,7'd33}:		p = 14'd1782;
            {7'd54,7'd34}:		p = 14'd1836;
            {7'd54,7'd35}:		p = 14'd1890;
            {7'd54,7'd36}:		p = 14'd1944;
            {7'd54,7'd37}:		p = 14'd1998;
            {7'd54,7'd38}:		p = 14'd2052;
            {7'd54,7'd39}:		p = 14'd2106;
            {7'd54,7'd40}:		p = 14'd2160;
            {7'd54,7'd41}:		p = 14'd2214;
            {7'd54,7'd42}:		p = 14'd2268;
            {7'd54,7'd43}:		p = 14'd2322;
            {7'd54,7'd44}:		p = 14'd2376;
            {7'd54,7'd45}:		p = 14'd2430;
            {7'd54,7'd46}:		p = 14'd2484;
            {7'd54,7'd47}:		p = 14'd2538;
            {7'd54,7'd48}:		p = 14'd2592;
            {7'd54,7'd49}:		p = 14'd2646;
            {7'd54,7'd50}:		p = 14'd2700;
            {7'd54,7'd51}:		p = 14'd2754;
            {7'd54,7'd52}:		p = 14'd2808;
            {7'd54,7'd53}:		p = 14'd2862;
            {7'd54,7'd54}:		p = 14'd2916;
            {7'd54,7'd55}:		p = 14'd2970;
            {7'd54,7'd56}:		p = 14'd3024;
            {7'd54,7'd57}:		p = 14'd3078;
            {7'd54,7'd58}:		p = 14'd3132;
            {7'd54,7'd59}:		p = 14'd3186;
            {7'd54,7'd60}:		p = 14'd3240;
            {7'd54,7'd61}:		p = 14'd3294;
            {7'd54,7'd62}:		p = 14'd3348;
            {7'd54,7'd63}:		p = 14'd3402;
            {7'd54,7'd64}:		p = 14'd3456;
            {7'd54,7'd65}:		p = 14'd3510;
            {7'd54,7'd66}:		p = 14'd3564;
            {7'd54,7'd67}:		p = 14'd3618;
            {7'd54,7'd68}:		p = 14'd3672;
            {7'd54,7'd69}:		p = 14'd3726;
            {7'd54,7'd70}:		p = 14'd3780;
            {7'd54,7'd71}:		p = 14'd3834;
            {7'd54,7'd72}:		p = 14'd3888;
            {7'd54,7'd73}:		p = 14'd3942;
            {7'd54,7'd74}:		p = 14'd3996;
            {7'd54,7'd75}:		p = 14'd4050;
            {7'd54,7'd76}:		p = 14'd4104;
            {7'd54,7'd77}:		p = 14'd4158;
            {7'd54,7'd78}:		p = 14'd4212;
            {7'd54,7'd79}:		p = 14'd4266;
            {7'd54,7'd80}:		p = 14'd4320;
            {7'd54,7'd81}:		p = 14'd4374;
            {7'd54,7'd82}:		p = 14'd4428;
            {7'd54,7'd83}:		p = 14'd4482;
            {7'd54,7'd84}:		p = 14'd4536;
            {7'd54,7'd85}:		p = 14'd4590;
            {7'd54,7'd86}:		p = 14'd4644;
            {7'd54,7'd87}:		p = 14'd4698;
            {7'd54,7'd88}:		p = 14'd4752;
            {7'd54,7'd89}:		p = 14'd4806;
            {7'd54,7'd90}:		p = 14'd4860;
            {7'd54,7'd91}:		p = 14'd4914;
            {7'd54,7'd92}:		p = 14'd4968;
            {7'd54,7'd93}:		p = 14'd5022;
            {7'd54,7'd94}:		p = 14'd5076;
            {7'd54,7'd95}:		p = 14'd5130;
            {7'd54,7'd96}:		p = 14'd5184;
            {7'd54,7'd97}:		p = 14'd5238;
            {7'd54,7'd98}:		p = 14'd5292;
            {7'd54,7'd99}:		p = 14'd5346;
            {7'd54,7'd100}:		p = 14'd5400;
            {7'd54,7'd101}:		p = 14'd5454;
            {7'd54,7'd102}:		p = 14'd5508;
            {7'd54,7'd103}:		p = 14'd5562;
            {7'd54,7'd104}:		p = 14'd5616;
            {7'd54,7'd105}:		p = 14'd5670;
            {7'd54,7'd106}:		p = 14'd5724;
            {7'd54,7'd107}:		p = 14'd5778;
            {7'd54,7'd108}:		p = 14'd5832;
            {7'd54,7'd109}:		p = 14'd5886;
            {7'd54,7'd110}:		p = 14'd5940;
            {7'd54,7'd111}:		p = 14'd5994;
            {7'd54,7'd112}:		p = 14'd6048;
            {7'd54,7'd113}:		p = 14'd6102;
            {7'd54,7'd114}:		p = 14'd6156;
            {7'd54,7'd115}:		p = 14'd6210;
            {7'd54,7'd116}:		p = 14'd6264;
            {7'd54,7'd117}:		p = 14'd6318;
            {7'd54,7'd118}:		p = 14'd6372;
            {7'd54,7'd119}:		p = 14'd6426;
            {7'd54,7'd120}:		p = 14'd6480;
            {7'd54,7'd121}:		p = 14'd6534;
            {7'd54,7'd122}:		p = 14'd6588;
            {7'd54,7'd123}:		p = 14'd6642;
            {7'd54,7'd124}:		p = 14'd6696;
            {7'd54,7'd125}:		p = 14'd6750;
            {7'd54,7'd126}:		p = 14'd6804;
            {7'd54,7'd127}:		p = 14'd6858;
            {7'd55,7'd0}:		p = 14'd0;
            {7'd55,7'd1}:		p = 14'd55;
            {7'd55,7'd2}:		p = 14'd110;
            {7'd55,7'd3}:		p = 14'd165;
            {7'd55,7'd4}:		p = 14'd220;
            {7'd55,7'd5}:		p = 14'd275;
            {7'd55,7'd6}:		p = 14'd330;
            {7'd55,7'd7}:		p = 14'd385;
            {7'd55,7'd8}:		p = 14'd440;
            {7'd55,7'd9}:		p = 14'd495;
            {7'd55,7'd10}:		p = 14'd550;
            {7'd55,7'd11}:		p = 14'd605;
            {7'd55,7'd12}:		p = 14'd660;
            {7'd55,7'd13}:		p = 14'd715;
            {7'd55,7'd14}:		p = 14'd770;
            {7'd55,7'd15}:		p = 14'd825;
            {7'd55,7'd16}:		p = 14'd880;
            {7'd55,7'd17}:		p = 14'd935;
            {7'd55,7'd18}:		p = 14'd990;
            {7'd55,7'd19}:		p = 14'd1045;
            {7'd55,7'd20}:		p = 14'd1100;
            {7'd55,7'd21}:		p = 14'd1155;
            {7'd55,7'd22}:		p = 14'd1210;
            {7'd55,7'd23}:		p = 14'd1265;
            {7'd55,7'd24}:		p = 14'd1320;
            {7'd55,7'd25}:		p = 14'd1375;
            {7'd55,7'd26}:		p = 14'd1430;
            {7'd55,7'd27}:		p = 14'd1485;
            {7'd55,7'd28}:		p = 14'd1540;
            {7'd55,7'd29}:		p = 14'd1595;
            {7'd55,7'd30}:		p = 14'd1650;
            {7'd55,7'd31}:		p = 14'd1705;
            {7'd55,7'd32}:		p = 14'd1760;
            {7'd55,7'd33}:		p = 14'd1815;
            {7'd55,7'd34}:		p = 14'd1870;
            {7'd55,7'd35}:		p = 14'd1925;
            {7'd55,7'd36}:		p = 14'd1980;
            {7'd55,7'd37}:		p = 14'd2035;
            {7'd55,7'd38}:		p = 14'd2090;
            {7'd55,7'd39}:		p = 14'd2145;
            {7'd55,7'd40}:		p = 14'd2200;
            {7'd55,7'd41}:		p = 14'd2255;
            {7'd55,7'd42}:		p = 14'd2310;
            {7'd55,7'd43}:		p = 14'd2365;
            {7'd55,7'd44}:		p = 14'd2420;
            {7'd55,7'd45}:		p = 14'd2475;
            {7'd55,7'd46}:		p = 14'd2530;
            {7'd55,7'd47}:		p = 14'd2585;
            {7'd55,7'd48}:		p = 14'd2640;
            {7'd55,7'd49}:		p = 14'd2695;
            {7'd55,7'd50}:		p = 14'd2750;
            {7'd55,7'd51}:		p = 14'd2805;
            {7'd55,7'd52}:		p = 14'd2860;
            {7'd55,7'd53}:		p = 14'd2915;
            {7'd55,7'd54}:		p = 14'd2970;
            {7'd55,7'd55}:		p = 14'd3025;
            {7'd55,7'd56}:		p = 14'd3080;
            {7'd55,7'd57}:		p = 14'd3135;
            {7'd55,7'd58}:		p = 14'd3190;
            {7'd55,7'd59}:		p = 14'd3245;
            {7'd55,7'd60}:		p = 14'd3300;
            {7'd55,7'd61}:		p = 14'd3355;
            {7'd55,7'd62}:		p = 14'd3410;
            {7'd55,7'd63}:		p = 14'd3465;
            {7'd55,7'd64}:		p = 14'd3520;
            {7'd55,7'd65}:		p = 14'd3575;
            {7'd55,7'd66}:		p = 14'd3630;
            {7'd55,7'd67}:		p = 14'd3685;
            {7'd55,7'd68}:		p = 14'd3740;
            {7'd55,7'd69}:		p = 14'd3795;
            {7'd55,7'd70}:		p = 14'd3850;
            {7'd55,7'd71}:		p = 14'd3905;
            {7'd55,7'd72}:		p = 14'd3960;
            {7'd55,7'd73}:		p = 14'd4015;
            {7'd55,7'd74}:		p = 14'd4070;
            {7'd55,7'd75}:		p = 14'd4125;
            {7'd55,7'd76}:		p = 14'd4180;
            {7'd55,7'd77}:		p = 14'd4235;
            {7'd55,7'd78}:		p = 14'd4290;
            {7'd55,7'd79}:		p = 14'd4345;
            {7'd55,7'd80}:		p = 14'd4400;
            {7'd55,7'd81}:		p = 14'd4455;
            {7'd55,7'd82}:		p = 14'd4510;
            {7'd55,7'd83}:		p = 14'd4565;
            {7'd55,7'd84}:		p = 14'd4620;
            {7'd55,7'd85}:		p = 14'd4675;
            {7'd55,7'd86}:		p = 14'd4730;
            {7'd55,7'd87}:		p = 14'd4785;
            {7'd55,7'd88}:		p = 14'd4840;
            {7'd55,7'd89}:		p = 14'd4895;
            {7'd55,7'd90}:		p = 14'd4950;
            {7'd55,7'd91}:		p = 14'd5005;
            {7'd55,7'd92}:		p = 14'd5060;
            {7'd55,7'd93}:		p = 14'd5115;
            {7'd55,7'd94}:		p = 14'd5170;
            {7'd55,7'd95}:		p = 14'd5225;
            {7'd55,7'd96}:		p = 14'd5280;
            {7'd55,7'd97}:		p = 14'd5335;
            {7'd55,7'd98}:		p = 14'd5390;
            {7'd55,7'd99}:		p = 14'd5445;
            {7'd55,7'd100}:		p = 14'd5500;
            {7'd55,7'd101}:		p = 14'd5555;
            {7'd55,7'd102}:		p = 14'd5610;
            {7'd55,7'd103}:		p = 14'd5665;
            {7'd55,7'd104}:		p = 14'd5720;
            {7'd55,7'd105}:		p = 14'd5775;
            {7'd55,7'd106}:		p = 14'd5830;
            {7'd55,7'd107}:		p = 14'd5885;
            {7'd55,7'd108}:		p = 14'd5940;
            {7'd55,7'd109}:		p = 14'd5995;
            {7'd55,7'd110}:		p = 14'd6050;
            {7'd55,7'd111}:		p = 14'd6105;
            {7'd55,7'd112}:		p = 14'd6160;
            {7'd55,7'd113}:		p = 14'd6215;
            {7'd55,7'd114}:		p = 14'd6270;
            {7'd55,7'd115}:		p = 14'd6325;
            {7'd55,7'd116}:		p = 14'd6380;
            {7'd55,7'd117}:		p = 14'd6435;
            {7'd55,7'd118}:		p = 14'd6490;
            {7'd55,7'd119}:		p = 14'd6545;
            {7'd55,7'd120}:		p = 14'd6600;
            {7'd55,7'd121}:		p = 14'd6655;
            {7'd55,7'd122}:		p = 14'd6710;
            {7'd55,7'd123}:		p = 14'd6765;
            {7'd55,7'd124}:		p = 14'd6820;
            {7'd55,7'd125}:		p = 14'd6875;
            {7'd55,7'd126}:		p = 14'd6930;
            {7'd55,7'd127}:		p = 14'd6985;
            {7'd56,7'd0}:		p = 14'd0;
            {7'd56,7'd1}:		p = 14'd56;
            {7'd56,7'd2}:		p = 14'd112;
            {7'd56,7'd3}:		p = 14'd168;
            {7'd56,7'd4}:		p = 14'd224;
            {7'd56,7'd5}:		p = 14'd280;
            {7'd56,7'd6}:		p = 14'd336;
            {7'd56,7'd7}:		p = 14'd392;
            {7'd56,7'd8}:		p = 14'd448;
            {7'd56,7'd9}:		p = 14'd504;
            {7'd56,7'd10}:		p = 14'd560;
            {7'd56,7'd11}:		p = 14'd616;
            {7'd56,7'd12}:		p = 14'd672;
            {7'd56,7'd13}:		p = 14'd728;
            {7'd56,7'd14}:		p = 14'd784;
            {7'd56,7'd15}:		p = 14'd840;
            {7'd56,7'd16}:		p = 14'd896;
            {7'd56,7'd17}:		p = 14'd952;
            {7'd56,7'd18}:		p = 14'd1008;
            {7'd56,7'd19}:		p = 14'd1064;
            {7'd56,7'd20}:		p = 14'd1120;
            {7'd56,7'd21}:		p = 14'd1176;
            {7'd56,7'd22}:		p = 14'd1232;
            {7'd56,7'd23}:		p = 14'd1288;
            {7'd56,7'd24}:		p = 14'd1344;
            {7'd56,7'd25}:		p = 14'd1400;
            {7'd56,7'd26}:		p = 14'd1456;
            {7'd56,7'd27}:		p = 14'd1512;
            {7'd56,7'd28}:		p = 14'd1568;
            {7'd56,7'd29}:		p = 14'd1624;
            {7'd56,7'd30}:		p = 14'd1680;
            {7'd56,7'd31}:		p = 14'd1736;
            {7'd56,7'd32}:		p = 14'd1792;
            {7'd56,7'd33}:		p = 14'd1848;
            {7'd56,7'd34}:		p = 14'd1904;
            {7'd56,7'd35}:		p = 14'd1960;
            {7'd56,7'd36}:		p = 14'd2016;
            {7'd56,7'd37}:		p = 14'd2072;
            {7'd56,7'd38}:		p = 14'd2128;
            {7'd56,7'd39}:		p = 14'd2184;
            {7'd56,7'd40}:		p = 14'd2240;
            {7'd56,7'd41}:		p = 14'd2296;
            {7'd56,7'd42}:		p = 14'd2352;
            {7'd56,7'd43}:		p = 14'd2408;
            {7'd56,7'd44}:		p = 14'd2464;
            {7'd56,7'd45}:		p = 14'd2520;
            {7'd56,7'd46}:		p = 14'd2576;
            {7'd56,7'd47}:		p = 14'd2632;
            {7'd56,7'd48}:		p = 14'd2688;
            {7'd56,7'd49}:		p = 14'd2744;
            {7'd56,7'd50}:		p = 14'd2800;
            {7'd56,7'd51}:		p = 14'd2856;
            {7'd56,7'd52}:		p = 14'd2912;
            {7'd56,7'd53}:		p = 14'd2968;
            {7'd56,7'd54}:		p = 14'd3024;
            {7'd56,7'd55}:		p = 14'd3080;
            {7'd56,7'd56}:		p = 14'd3136;
            {7'd56,7'd57}:		p = 14'd3192;
            {7'd56,7'd58}:		p = 14'd3248;
            {7'd56,7'd59}:		p = 14'd3304;
            {7'd56,7'd60}:		p = 14'd3360;
            {7'd56,7'd61}:		p = 14'd3416;
            {7'd56,7'd62}:		p = 14'd3472;
            {7'd56,7'd63}:		p = 14'd3528;
            {7'd56,7'd64}:		p = 14'd3584;
            {7'd56,7'd65}:		p = 14'd3640;
            {7'd56,7'd66}:		p = 14'd3696;
            {7'd56,7'd67}:		p = 14'd3752;
            {7'd56,7'd68}:		p = 14'd3808;
            {7'd56,7'd69}:		p = 14'd3864;
            {7'd56,7'd70}:		p = 14'd3920;
            {7'd56,7'd71}:		p = 14'd3976;
            {7'd56,7'd72}:		p = 14'd4032;
            {7'd56,7'd73}:		p = 14'd4088;
            {7'd56,7'd74}:		p = 14'd4144;
            {7'd56,7'd75}:		p = 14'd4200;
            {7'd56,7'd76}:		p = 14'd4256;
            {7'd56,7'd77}:		p = 14'd4312;
            {7'd56,7'd78}:		p = 14'd4368;
            {7'd56,7'd79}:		p = 14'd4424;
            {7'd56,7'd80}:		p = 14'd4480;
            {7'd56,7'd81}:		p = 14'd4536;
            {7'd56,7'd82}:		p = 14'd4592;
            {7'd56,7'd83}:		p = 14'd4648;
            {7'd56,7'd84}:		p = 14'd4704;
            {7'd56,7'd85}:		p = 14'd4760;
            {7'd56,7'd86}:		p = 14'd4816;
            {7'd56,7'd87}:		p = 14'd4872;
            {7'd56,7'd88}:		p = 14'd4928;
            {7'd56,7'd89}:		p = 14'd4984;
            {7'd56,7'd90}:		p = 14'd5040;
            {7'd56,7'd91}:		p = 14'd5096;
            {7'd56,7'd92}:		p = 14'd5152;
            {7'd56,7'd93}:		p = 14'd5208;
            {7'd56,7'd94}:		p = 14'd5264;
            {7'd56,7'd95}:		p = 14'd5320;
            {7'd56,7'd96}:		p = 14'd5376;
            {7'd56,7'd97}:		p = 14'd5432;
            {7'd56,7'd98}:		p = 14'd5488;
            {7'd56,7'd99}:		p = 14'd5544;
            {7'd56,7'd100}:		p = 14'd5600;
            {7'd56,7'd101}:		p = 14'd5656;
            {7'd56,7'd102}:		p = 14'd5712;
            {7'd56,7'd103}:		p = 14'd5768;
            {7'd56,7'd104}:		p = 14'd5824;
            {7'd56,7'd105}:		p = 14'd5880;
            {7'd56,7'd106}:		p = 14'd5936;
            {7'd56,7'd107}:		p = 14'd5992;
            {7'd56,7'd108}:		p = 14'd6048;
            {7'd56,7'd109}:		p = 14'd6104;
            {7'd56,7'd110}:		p = 14'd6160;
            {7'd56,7'd111}:		p = 14'd6216;
            {7'd56,7'd112}:		p = 14'd6272;
            {7'd56,7'd113}:		p = 14'd6328;
            {7'd56,7'd114}:		p = 14'd6384;
            {7'd56,7'd115}:		p = 14'd6440;
            {7'd56,7'd116}:		p = 14'd6496;
            {7'd56,7'd117}:		p = 14'd6552;
            {7'd56,7'd118}:		p = 14'd6608;
            {7'd56,7'd119}:		p = 14'd6664;
            {7'd56,7'd120}:		p = 14'd6720;
            {7'd56,7'd121}:		p = 14'd6776;
            {7'd56,7'd122}:		p = 14'd6832;
            {7'd56,7'd123}:		p = 14'd6888;
            {7'd56,7'd124}:		p = 14'd6944;
            {7'd56,7'd125}:		p = 14'd7000;
            {7'd56,7'd126}:		p = 14'd7056;
            {7'd56,7'd127}:		p = 14'd7112;
            {7'd57,7'd0}:		p = 14'd0;
            {7'd57,7'd1}:		p = 14'd57;
            {7'd57,7'd2}:		p = 14'd114;
            {7'd57,7'd3}:		p = 14'd171;
            {7'd57,7'd4}:		p = 14'd228;
            {7'd57,7'd5}:		p = 14'd285;
            {7'd57,7'd6}:		p = 14'd342;
            {7'd57,7'd7}:		p = 14'd399;
            {7'd57,7'd8}:		p = 14'd456;
            {7'd57,7'd9}:		p = 14'd513;
            {7'd57,7'd10}:		p = 14'd570;
            {7'd57,7'd11}:		p = 14'd627;
            {7'd57,7'd12}:		p = 14'd684;
            {7'd57,7'd13}:		p = 14'd741;
            {7'd57,7'd14}:		p = 14'd798;
            {7'd57,7'd15}:		p = 14'd855;
            {7'd57,7'd16}:		p = 14'd912;
            {7'd57,7'd17}:		p = 14'd969;
            {7'd57,7'd18}:		p = 14'd1026;
            {7'd57,7'd19}:		p = 14'd1083;
            {7'd57,7'd20}:		p = 14'd1140;
            {7'd57,7'd21}:		p = 14'd1197;
            {7'd57,7'd22}:		p = 14'd1254;
            {7'd57,7'd23}:		p = 14'd1311;
            {7'd57,7'd24}:		p = 14'd1368;
            {7'd57,7'd25}:		p = 14'd1425;
            {7'd57,7'd26}:		p = 14'd1482;
            {7'd57,7'd27}:		p = 14'd1539;
            {7'd57,7'd28}:		p = 14'd1596;
            {7'd57,7'd29}:		p = 14'd1653;
            {7'd57,7'd30}:		p = 14'd1710;
            {7'd57,7'd31}:		p = 14'd1767;
            {7'd57,7'd32}:		p = 14'd1824;
            {7'd57,7'd33}:		p = 14'd1881;
            {7'd57,7'd34}:		p = 14'd1938;
            {7'd57,7'd35}:		p = 14'd1995;
            {7'd57,7'd36}:		p = 14'd2052;
            {7'd57,7'd37}:		p = 14'd2109;
            {7'd57,7'd38}:		p = 14'd2166;
            {7'd57,7'd39}:		p = 14'd2223;
            {7'd57,7'd40}:		p = 14'd2280;
            {7'd57,7'd41}:		p = 14'd2337;
            {7'd57,7'd42}:		p = 14'd2394;
            {7'd57,7'd43}:		p = 14'd2451;
            {7'd57,7'd44}:		p = 14'd2508;
            {7'd57,7'd45}:		p = 14'd2565;
            {7'd57,7'd46}:		p = 14'd2622;
            {7'd57,7'd47}:		p = 14'd2679;
            {7'd57,7'd48}:		p = 14'd2736;
            {7'd57,7'd49}:		p = 14'd2793;
            {7'd57,7'd50}:		p = 14'd2850;
            {7'd57,7'd51}:		p = 14'd2907;
            {7'd57,7'd52}:		p = 14'd2964;
            {7'd57,7'd53}:		p = 14'd3021;
            {7'd57,7'd54}:		p = 14'd3078;
            {7'd57,7'd55}:		p = 14'd3135;
            {7'd57,7'd56}:		p = 14'd3192;
            {7'd57,7'd57}:		p = 14'd3249;
            {7'd57,7'd58}:		p = 14'd3306;
            {7'd57,7'd59}:		p = 14'd3363;
            {7'd57,7'd60}:		p = 14'd3420;
            {7'd57,7'd61}:		p = 14'd3477;
            {7'd57,7'd62}:		p = 14'd3534;
            {7'd57,7'd63}:		p = 14'd3591;
            {7'd57,7'd64}:		p = 14'd3648;
            {7'd57,7'd65}:		p = 14'd3705;
            {7'd57,7'd66}:		p = 14'd3762;
            {7'd57,7'd67}:		p = 14'd3819;
            {7'd57,7'd68}:		p = 14'd3876;
            {7'd57,7'd69}:		p = 14'd3933;
            {7'd57,7'd70}:		p = 14'd3990;
            {7'd57,7'd71}:		p = 14'd4047;
            {7'd57,7'd72}:		p = 14'd4104;
            {7'd57,7'd73}:		p = 14'd4161;
            {7'd57,7'd74}:		p = 14'd4218;
            {7'd57,7'd75}:		p = 14'd4275;
            {7'd57,7'd76}:		p = 14'd4332;
            {7'd57,7'd77}:		p = 14'd4389;
            {7'd57,7'd78}:		p = 14'd4446;
            {7'd57,7'd79}:		p = 14'd4503;
            {7'd57,7'd80}:		p = 14'd4560;
            {7'd57,7'd81}:		p = 14'd4617;
            {7'd57,7'd82}:		p = 14'd4674;
            {7'd57,7'd83}:		p = 14'd4731;
            {7'd57,7'd84}:		p = 14'd4788;
            {7'd57,7'd85}:		p = 14'd4845;
            {7'd57,7'd86}:		p = 14'd4902;
            {7'd57,7'd87}:		p = 14'd4959;
            {7'd57,7'd88}:		p = 14'd5016;
            {7'd57,7'd89}:		p = 14'd5073;
            {7'd57,7'd90}:		p = 14'd5130;
            {7'd57,7'd91}:		p = 14'd5187;
            {7'd57,7'd92}:		p = 14'd5244;
            {7'd57,7'd93}:		p = 14'd5301;
            {7'd57,7'd94}:		p = 14'd5358;
            {7'd57,7'd95}:		p = 14'd5415;
            {7'd57,7'd96}:		p = 14'd5472;
            {7'd57,7'd97}:		p = 14'd5529;
            {7'd57,7'd98}:		p = 14'd5586;
            {7'd57,7'd99}:		p = 14'd5643;
            {7'd57,7'd100}:		p = 14'd5700;
            {7'd57,7'd101}:		p = 14'd5757;
            {7'd57,7'd102}:		p = 14'd5814;
            {7'd57,7'd103}:		p = 14'd5871;
            {7'd57,7'd104}:		p = 14'd5928;
            {7'd57,7'd105}:		p = 14'd5985;
            {7'd57,7'd106}:		p = 14'd6042;
            {7'd57,7'd107}:		p = 14'd6099;
            {7'd57,7'd108}:		p = 14'd6156;
            {7'd57,7'd109}:		p = 14'd6213;
            {7'd57,7'd110}:		p = 14'd6270;
            {7'd57,7'd111}:		p = 14'd6327;
            {7'd57,7'd112}:		p = 14'd6384;
            {7'd57,7'd113}:		p = 14'd6441;
            {7'd57,7'd114}:		p = 14'd6498;
            {7'd57,7'd115}:		p = 14'd6555;
            {7'd57,7'd116}:		p = 14'd6612;
            {7'd57,7'd117}:		p = 14'd6669;
            {7'd57,7'd118}:		p = 14'd6726;
            {7'd57,7'd119}:		p = 14'd6783;
            {7'd57,7'd120}:		p = 14'd6840;
            {7'd57,7'd121}:		p = 14'd6897;
            {7'd57,7'd122}:		p = 14'd6954;
            {7'd57,7'd123}:		p = 14'd7011;
            {7'd57,7'd124}:		p = 14'd7068;
            {7'd57,7'd125}:		p = 14'd7125;
            {7'd57,7'd126}:		p = 14'd7182;
            {7'd57,7'd127}:		p = 14'd7239;
            {7'd58,7'd0}:		p = 14'd0;
            {7'd58,7'd1}:		p = 14'd58;
            {7'd58,7'd2}:		p = 14'd116;
            {7'd58,7'd3}:		p = 14'd174;
            {7'd58,7'd4}:		p = 14'd232;
            {7'd58,7'd5}:		p = 14'd290;
            {7'd58,7'd6}:		p = 14'd348;
            {7'd58,7'd7}:		p = 14'd406;
            {7'd58,7'd8}:		p = 14'd464;
            {7'd58,7'd9}:		p = 14'd522;
            {7'd58,7'd10}:		p = 14'd580;
            {7'd58,7'd11}:		p = 14'd638;
            {7'd58,7'd12}:		p = 14'd696;
            {7'd58,7'd13}:		p = 14'd754;
            {7'd58,7'd14}:		p = 14'd812;
            {7'd58,7'd15}:		p = 14'd870;
            {7'd58,7'd16}:		p = 14'd928;
            {7'd58,7'd17}:		p = 14'd986;
            {7'd58,7'd18}:		p = 14'd1044;
            {7'd58,7'd19}:		p = 14'd1102;
            {7'd58,7'd20}:		p = 14'd1160;
            {7'd58,7'd21}:		p = 14'd1218;
            {7'd58,7'd22}:		p = 14'd1276;
            {7'd58,7'd23}:		p = 14'd1334;
            {7'd58,7'd24}:		p = 14'd1392;
            {7'd58,7'd25}:		p = 14'd1450;
            {7'd58,7'd26}:		p = 14'd1508;
            {7'd58,7'd27}:		p = 14'd1566;
            {7'd58,7'd28}:		p = 14'd1624;
            {7'd58,7'd29}:		p = 14'd1682;
            {7'd58,7'd30}:		p = 14'd1740;
            {7'd58,7'd31}:		p = 14'd1798;
            {7'd58,7'd32}:		p = 14'd1856;
            {7'd58,7'd33}:		p = 14'd1914;
            {7'd58,7'd34}:		p = 14'd1972;
            {7'd58,7'd35}:		p = 14'd2030;
            {7'd58,7'd36}:		p = 14'd2088;
            {7'd58,7'd37}:		p = 14'd2146;
            {7'd58,7'd38}:		p = 14'd2204;
            {7'd58,7'd39}:		p = 14'd2262;
            {7'd58,7'd40}:		p = 14'd2320;
            {7'd58,7'd41}:		p = 14'd2378;
            {7'd58,7'd42}:		p = 14'd2436;
            {7'd58,7'd43}:		p = 14'd2494;
            {7'd58,7'd44}:		p = 14'd2552;
            {7'd58,7'd45}:		p = 14'd2610;
            {7'd58,7'd46}:		p = 14'd2668;
            {7'd58,7'd47}:		p = 14'd2726;
            {7'd58,7'd48}:		p = 14'd2784;
            {7'd58,7'd49}:		p = 14'd2842;
            {7'd58,7'd50}:		p = 14'd2900;
            {7'd58,7'd51}:		p = 14'd2958;
            {7'd58,7'd52}:		p = 14'd3016;
            {7'd58,7'd53}:		p = 14'd3074;
            {7'd58,7'd54}:		p = 14'd3132;
            {7'd58,7'd55}:		p = 14'd3190;
            {7'd58,7'd56}:		p = 14'd3248;
            {7'd58,7'd57}:		p = 14'd3306;
            {7'd58,7'd58}:		p = 14'd3364;
            {7'd58,7'd59}:		p = 14'd3422;
            {7'd58,7'd60}:		p = 14'd3480;
            {7'd58,7'd61}:		p = 14'd3538;
            {7'd58,7'd62}:		p = 14'd3596;
            {7'd58,7'd63}:		p = 14'd3654;
            {7'd58,7'd64}:		p = 14'd3712;
            {7'd58,7'd65}:		p = 14'd3770;
            {7'd58,7'd66}:		p = 14'd3828;
            {7'd58,7'd67}:		p = 14'd3886;
            {7'd58,7'd68}:		p = 14'd3944;
            {7'd58,7'd69}:		p = 14'd4002;
            {7'd58,7'd70}:		p = 14'd4060;
            {7'd58,7'd71}:		p = 14'd4118;
            {7'd58,7'd72}:		p = 14'd4176;
            {7'd58,7'd73}:		p = 14'd4234;
            {7'd58,7'd74}:		p = 14'd4292;
            {7'd58,7'd75}:		p = 14'd4350;
            {7'd58,7'd76}:		p = 14'd4408;
            {7'd58,7'd77}:		p = 14'd4466;
            {7'd58,7'd78}:		p = 14'd4524;
            {7'd58,7'd79}:		p = 14'd4582;
            {7'd58,7'd80}:		p = 14'd4640;
            {7'd58,7'd81}:		p = 14'd4698;
            {7'd58,7'd82}:		p = 14'd4756;
            {7'd58,7'd83}:		p = 14'd4814;
            {7'd58,7'd84}:		p = 14'd4872;
            {7'd58,7'd85}:		p = 14'd4930;
            {7'd58,7'd86}:		p = 14'd4988;
            {7'd58,7'd87}:		p = 14'd5046;
            {7'd58,7'd88}:		p = 14'd5104;
            {7'd58,7'd89}:		p = 14'd5162;
            {7'd58,7'd90}:		p = 14'd5220;
            {7'd58,7'd91}:		p = 14'd5278;
            {7'd58,7'd92}:		p = 14'd5336;
            {7'd58,7'd93}:		p = 14'd5394;
            {7'd58,7'd94}:		p = 14'd5452;
            {7'd58,7'd95}:		p = 14'd5510;
            {7'd58,7'd96}:		p = 14'd5568;
            {7'd58,7'd97}:		p = 14'd5626;
            {7'd58,7'd98}:		p = 14'd5684;
            {7'd58,7'd99}:		p = 14'd5742;
            {7'd58,7'd100}:		p = 14'd5800;
            {7'd58,7'd101}:		p = 14'd5858;
            {7'd58,7'd102}:		p = 14'd5916;
            {7'd58,7'd103}:		p = 14'd5974;
            {7'd58,7'd104}:		p = 14'd6032;
            {7'd58,7'd105}:		p = 14'd6090;
            {7'd58,7'd106}:		p = 14'd6148;
            {7'd58,7'd107}:		p = 14'd6206;
            {7'd58,7'd108}:		p = 14'd6264;
            {7'd58,7'd109}:		p = 14'd6322;
            {7'd58,7'd110}:		p = 14'd6380;
            {7'd58,7'd111}:		p = 14'd6438;
            {7'd58,7'd112}:		p = 14'd6496;
            {7'd58,7'd113}:		p = 14'd6554;
            {7'd58,7'd114}:		p = 14'd6612;
            {7'd58,7'd115}:		p = 14'd6670;
            {7'd58,7'd116}:		p = 14'd6728;
            {7'd58,7'd117}:		p = 14'd6786;
            {7'd58,7'd118}:		p = 14'd6844;
            {7'd58,7'd119}:		p = 14'd6902;
            {7'd58,7'd120}:		p = 14'd6960;
            {7'd58,7'd121}:		p = 14'd7018;
            {7'd58,7'd122}:		p = 14'd7076;
            {7'd58,7'd123}:		p = 14'd7134;
            {7'd58,7'd124}:		p = 14'd7192;
            {7'd58,7'd125}:		p = 14'd7250;
            {7'd58,7'd126}:		p = 14'd7308;
            {7'd58,7'd127}:		p = 14'd7366;
            {7'd59,7'd0}:		p = 14'd0;
            {7'd59,7'd1}:		p = 14'd59;
            {7'd59,7'd2}:		p = 14'd118;
            {7'd59,7'd3}:		p = 14'd177;
            {7'd59,7'd4}:		p = 14'd236;
            {7'd59,7'd5}:		p = 14'd295;
            {7'd59,7'd6}:		p = 14'd354;
            {7'd59,7'd7}:		p = 14'd413;
            {7'd59,7'd8}:		p = 14'd472;
            {7'd59,7'd9}:		p = 14'd531;
            {7'd59,7'd10}:		p = 14'd590;
            {7'd59,7'd11}:		p = 14'd649;
            {7'd59,7'd12}:		p = 14'd708;
            {7'd59,7'd13}:		p = 14'd767;
            {7'd59,7'd14}:		p = 14'd826;
            {7'd59,7'd15}:		p = 14'd885;
            {7'd59,7'd16}:		p = 14'd944;
            {7'd59,7'd17}:		p = 14'd1003;
            {7'd59,7'd18}:		p = 14'd1062;
            {7'd59,7'd19}:		p = 14'd1121;
            {7'd59,7'd20}:		p = 14'd1180;
            {7'd59,7'd21}:		p = 14'd1239;
            {7'd59,7'd22}:		p = 14'd1298;
            {7'd59,7'd23}:		p = 14'd1357;
            {7'd59,7'd24}:		p = 14'd1416;
            {7'd59,7'd25}:		p = 14'd1475;
            {7'd59,7'd26}:		p = 14'd1534;
            {7'd59,7'd27}:		p = 14'd1593;
            {7'd59,7'd28}:		p = 14'd1652;
            {7'd59,7'd29}:		p = 14'd1711;
            {7'd59,7'd30}:		p = 14'd1770;
            {7'd59,7'd31}:		p = 14'd1829;
            {7'd59,7'd32}:		p = 14'd1888;
            {7'd59,7'd33}:		p = 14'd1947;
            {7'd59,7'd34}:		p = 14'd2006;
            {7'd59,7'd35}:		p = 14'd2065;
            {7'd59,7'd36}:		p = 14'd2124;
            {7'd59,7'd37}:		p = 14'd2183;
            {7'd59,7'd38}:		p = 14'd2242;
            {7'd59,7'd39}:		p = 14'd2301;
            {7'd59,7'd40}:		p = 14'd2360;
            {7'd59,7'd41}:		p = 14'd2419;
            {7'd59,7'd42}:		p = 14'd2478;
            {7'd59,7'd43}:		p = 14'd2537;
            {7'd59,7'd44}:		p = 14'd2596;
            {7'd59,7'd45}:		p = 14'd2655;
            {7'd59,7'd46}:		p = 14'd2714;
            {7'd59,7'd47}:		p = 14'd2773;
            {7'd59,7'd48}:		p = 14'd2832;
            {7'd59,7'd49}:		p = 14'd2891;
            {7'd59,7'd50}:		p = 14'd2950;
            {7'd59,7'd51}:		p = 14'd3009;
            {7'd59,7'd52}:		p = 14'd3068;
            {7'd59,7'd53}:		p = 14'd3127;
            {7'd59,7'd54}:		p = 14'd3186;
            {7'd59,7'd55}:		p = 14'd3245;
            {7'd59,7'd56}:		p = 14'd3304;
            {7'd59,7'd57}:		p = 14'd3363;
            {7'd59,7'd58}:		p = 14'd3422;
            {7'd59,7'd59}:		p = 14'd3481;
            {7'd59,7'd60}:		p = 14'd3540;
            {7'd59,7'd61}:		p = 14'd3599;
            {7'd59,7'd62}:		p = 14'd3658;
            {7'd59,7'd63}:		p = 14'd3717;
            {7'd59,7'd64}:		p = 14'd3776;
            {7'd59,7'd65}:		p = 14'd3835;
            {7'd59,7'd66}:		p = 14'd3894;
            {7'd59,7'd67}:		p = 14'd3953;
            {7'd59,7'd68}:		p = 14'd4012;
            {7'd59,7'd69}:		p = 14'd4071;
            {7'd59,7'd70}:		p = 14'd4130;
            {7'd59,7'd71}:		p = 14'd4189;
            {7'd59,7'd72}:		p = 14'd4248;
            {7'd59,7'd73}:		p = 14'd4307;
            {7'd59,7'd74}:		p = 14'd4366;
            {7'd59,7'd75}:		p = 14'd4425;
            {7'd59,7'd76}:		p = 14'd4484;
            {7'd59,7'd77}:		p = 14'd4543;
            {7'd59,7'd78}:		p = 14'd4602;
            {7'd59,7'd79}:		p = 14'd4661;
            {7'd59,7'd80}:		p = 14'd4720;
            {7'd59,7'd81}:		p = 14'd4779;
            {7'd59,7'd82}:		p = 14'd4838;
            {7'd59,7'd83}:		p = 14'd4897;
            {7'd59,7'd84}:		p = 14'd4956;
            {7'd59,7'd85}:		p = 14'd5015;
            {7'd59,7'd86}:		p = 14'd5074;
            {7'd59,7'd87}:		p = 14'd5133;
            {7'd59,7'd88}:		p = 14'd5192;
            {7'd59,7'd89}:		p = 14'd5251;
            {7'd59,7'd90}:		p = 14'd5310;
            {7'd59,7'd91}:		p = 14'd5369;
            {7'd59,7'd92}:		p = 14'd5428;
            {7'd59,7'd93}:		p = 14'd5487;
            {7'd59,7'd94}:		p = 14'd5546;
            {7'd59,7'd95}:		p = 14'd5605;
            {7'd59,7'd96}:		p = 14'd5664;
            {7'd59,7'd97}:		p = 14'd5723;
            {7'd59,7'd98}:		p = 14'd5782;
            {7'd59,7'd99}:		p = 14'd5841;
            {7'd59,7'd100}:		p = 14'd5900;
            {7'd59,7'd101}:		p = 14'd5959;
            {7'd59,7'd102}:		p = 14'd6018;
            {7'd59,7'd103}:		p = 14'd6077;
            {7'd59,7'd104}:		p = 14'd6136;
            {7'd59,7'd105}:		p = 14'd6195;
            {7'd59,7'd106}:		p = 14'd6254;
            {7'd59,7'd107}:		p = 14'd6313;
            {7'd59,7'd108}:		p = 14'd6372;
            {7'd59,7'd109}:		p = 14'd6431;
            {7'd59,7'd110}:		p = 14'd6490;
            {7'd59,7'd111}:		p = 14'd6549;
            {7'd59,7'd112}:		p = 14'd6608;
            {7'd59,7'd113}:		p = 14'd6667;
            {7'd59,7'd114}:		p = 14'd6726;
            {7'd59,7'd115}:		p = 14'd6785;
            {7'd59,7'd116}:		p = 14'd6844;
            {7'd59,7'd117}:		p = 14'd6903;
            {7'd59,7'd118}:		p = 14'd6962;
            {7'd59,7'd119}:		p = 14'd7021;
            {7'd59,7'd120}:		p = 14'd7080;
            {7'd59,7'd121}:		p = 14'd7139;
            {7'd59,7'd122}:		p = 14'd7198;
            {7'd59,7'd123}:		p = 14'd7257;
            {7'd59,7'd124}:		p = 14'd7316;
            {7'd59,7'd125}:		p = 14'd7375;
            {7'd59,7'd126}:		p = 14'd7434;
            {7'd59,7'd127}:		p = 14'd7493;
            {7'd60,7'd0}:		p = 14'd0;
            {7'd60,7'd1}:		p = 14'd60;
            {7'd60,7'd2}:		p = 14'd120;
            {7'd60,7'd3}:		p = 14'd180;
            {7'd60,7'd4}:		p = 14'd240;
            {7'd60,7'd5}:		p = 14'd300;
            {7'd60,7'd6}:		p = 14'd360;
            {7'd60,7'd7}:		p = 14'd420;
            {7'd60,7'd8}:		p = 14'd480;
            {7'd60,7'd9}:		p = 14'd540;
            {7'd60,7'd10}:		p = 14'd600;
            {7'd60,7'd11}:		p = 14'd660;
            {7'd60,7'd12}:		p = 14'd720;
            {7'd60,7'd13}:		p = 14'd780;
            {7'd60,7'd14}:		p = 14'd840;
            {7'd60,7'd15}:		p = 14'd900;
            {7'd60,7'd16}:		p = 14'd960;
            {7'd60,7'd17}:		p = 14'd1020;
            {7'd60,7'd18}:		p = 14'd1080;
            {7'd60,7'd19}:		p = 14'd1140;
            {7'd60,7'd20}:		p = 14'd1200;
            {7'd60,7'd21}:		p = 14'd1260;
            {7'd60,7'd22}:		p = 14'd1320;
            {7'd60,7'd23}:		p = 14'd1380;
            {7'd60,7'd24}:		p = 14'd1440;
            {7'd60,7'd25}:		p = 14'd1500;
            {7'd60,7'd26}:		p = 14'd1560;
            {7'd60,7'd27}:		p = 14'd1620;
            {7'd60,7'd28}:		p = 14'd1680;
            {7'd60,7'd29}:		p = 14'd1740;
            {7'd60,7'd30}:		p = 14'd1800;
            {7'd60,7'd31}:		p = 14'd1860;
            {7'd60,7'd32}:		p = 14'd1920;
            {7'd60,7'd33}:		p = 14'd1980;
            {7'd60,7'd34}:		p = 14'd2040;
            {7'd60,7'd35}:		p = 14'd2100;
            {7'd60,7'd36}:		p = 14'd2160;
            {7'd60,7'd37}:		p = 14'd2220;
            {7'd60,7'd38}:		p = 14'd2280;
            {7'd60,7'd39}:		p = 14'd2340;
            {7'd60,7'd40}:		p = 14'd2400;
            {7'd60,7'd41}:		p = 14'd2460;
            {7'd60,7'd42}:		p = 14'd2520;
            {7'd60,7'd43}:		p = 14'd2580;
            {7'd60,7'd44}:		p = 14'd2640;
            {7'd60,7'd45}:		p = 14'd2700;
            {7'd60,7'd46}:		p = 14'd2760;
            {7'd60,7'd47}:		p = 14'd2820;
            {7'd60,7'd48}:		p = 14'd2880;
            {7'd60,7'd49}:		p = 14'd2940;
            {7'd60,7'd50}:		p = 14'd3000;
            {7'd60,7'd51}:		p = 14'd3060;
            {7'd60,7'd52}:		p = 14'd3120;
            {7'd60,7'd53}:		p = 14'd3180;
            {7'd60,7'd54}:		p = 14'd3240;
            {7'd60,7'd55}:		p = 14'd3300;
            {7'd60,7'd56}:		p = 14'd3360;
            {7'd60,7'd57}:		p = 14'd3420;
            {7'd60,7'd58}:		p = 14'd3480;
            {7'd60,7'd59}:		p = 14'd3540;
            {7'd60,7'd60}:		p = 14'd3600;
            {7'd60,7'd61}:		p = 14'd3660;
            {7'd60,7'd62}:		p = 14'd3720;
            {7'd60,7'd63}:		p = 14'd3780;
            {7'd60,7'd64}:		p = 14'd3840;
            {7'd60,7'd65}:		p = 14'd3900;
            {7'd60,7'd66}:		p = 14'd3960;
            {7'd60,7'd67}:		p = 14'd4020;
            {7'd60,7'd68}:		p = 14'd4080;
            {7'd60,7'd69}:		p = 14'd4140;
            {7'd60,7'd70}:		p = 14'd4200;
            {7'd60,7'd71}:		p = 14'd4260;
            {7'd60,7'd72}:		p = 14'd4320;
            {7'd60,7'd73}:		p = 14'd4380;
            {7'd60,7'd74}:		p = 14'd4440;
            {7'd60,7'd75}:		p = 14'd4500;
            {7'd60,7'd76}:		p = 14'd4560;
            {7'd60,7'd77}:		p = 14'd4620;
            {7'd60,7'd78}:		p = 14'd4680;
            {7'd60,7'd79}:		p = 14'd4740;
            {7'd60,7'd80}:		p = 14'd4800;
            {7'd60,7'd81}:		p = 14'd4860;
            {7'd60,7'd82}:		p = 14'd4920;
            {7'd60,7'd83}:		p = 14'd4980;
            {7'd60,7'd84}:		p = 14'd5040;
            {7'd60,7'd85}:		p = 14'd5100;
            {7'd60,7'd86}:		p = 14'd5160;
            {7'd60,7'd87}:		p = 14'd5220;
            {7'd60,7'd88}:		p = 14'd5280;
            {7'd60,7'd89}:		p = 14'd5340;
            {7'd60,7'd90}:		p = 14'd5400;
            {7'd60,7'd91}:		p = 14'd5460;
            {7'd60,7'd92}:		p = 14'd5520;
            {7'd60,7'd93}:		p = 14'd5580;
            {7'd60,7'd94}:		p = 14'd5640;
            {7'd60,7'd95}:		p = 14'd5700;
            {7'd60,7'd96}:		p = 14'd5760;
            {7'd60,7'd97}:		p = 14'd5820;
            {7'd60,7'd98}:		p = 14'd5880;
            {7'd60,7'd99}:		p = 14'd5940;
            {7'd60,7'd100}:		p = 14'd6000;
            {7'd60,7'd101}:		p = 14'd6060;
            {7'd60,7'd102}:		p = 14'd6120;
            {7'd60,7'd103}:		p = 14'd6180;
            {7'd60,7'd104}:		p = 14'd6240;
            {7'd60,7'd105}:		p = 14'd6300;
            {7'd60,7'd106}:		p = 14'd6360;
            {7'd60,7'd107}:		p = 14'd6420;
            {7'd60,7'd108}:		p = 14'd6480;
            {7'd60,7'd109}:		p = 14'd6540;
            {7'd60,7'd110}:		p = 14'd6600;
            {7'd60,7'd111}:		p = 14'd6660;
            {7'd60,7'd112}:		p = 14'd6720;
            {7'd60,7'd113}:		p = 14'd6780;
            {7'd60,7'd114}:		p = 14'd6840;
            {7'd60,7'd115}:		p = 14'd6900;
            {7'd60,7'd116}:		p = 14'd6960;
            {7'd60,7'd117}:		p = 14'd7020;
            {7'd60,7'd118}:		p = 14'd7080;
            {7'd60,7'd119}:		p = 14'd7140;
            {7'd60,7'd120}:		p = 14'd7200;
            {7'd60,7'd121}:		p = 14'd7260;
            {7'd60,7'd122}:		p = 14'd7320;
            {7'd60,7'd123}:		p = 14'd7380;
            {7'd60,7'd124}:		p = 14'd7440;
            {7'd60,7'd125}:		p = 14'd7500;
            {7'd60,7'd126}:		p = 14'd7560;
            {7'd60,7'd127}:		p = 14'd7620;
            {7'd61,7'd0}:		p = 14'd0;
            {7'd61,7'd1}:		p = 14'd61;
            {7'd61,7'd2}:		p = 14'd122;
            {7'd61,7'd3}:		p = 14'd183;
            {7'd61,7'd4}:		p = 14'd244;
            {7'd61,7'd5}:		p = 14'd305;
            {7'd61,7'd6}:		p = 14'd366;
            {7'd61,7'd7}:		p = 14'd427;
            {7'd61,7'd8}:		p = 14'd488;
            {7'd61,7'd9}:		p = 14'd549;
            {7'd61,7'd10}:		p = 14'd610;
            {7'd61,7'd11}:		p = 14'd671;
            {7'd61,7'd12}:		p = 14'd732;
            {7'd61,7'd13}:		p = 14'd793;
            {7'd61,7'd14}:		p = 14'd854;
            {7'd61,7'd15}:		p = 14'd915;
            {7'd61,7'd16}:		p = 14'd976;
            {7'd61,7'd17}:		p = 14'd1037;
            {7'd61,7'd18}:		p = 14'd1098;
            {7'd61,7'd19}:		p = 14'd1159;
            {7'd61,7'd20}:		p = 14'd1220;
            {7'd61,7'd21}:		p = 14'd1281;
            {7'd61,7'd22}:		p = 14'd1342;
            {7'd61,7'd23}:		p = 14'd1403;
            {7'd61,7'd24}:		p = 14'd1464;
            {7'd61,7'd25}:		p = 14'd1525;
            {7'd61,7'd26}:		p = 14'd1586;
            {7'd61,7'd27}:		p = 14'd1647;
            {7'd61,7'd28}:		p = 14'd1708;
            {7'd61,7'd29}:		p = 14'd1769;
            {7'd61,7'd30}:		p = 14'd1830;
            {7'd61,7'd31}:		p = 14'd1891;
            {7'd61,7'd32}:		p = 14'd1952;
            {7'd61,7'd33}:		p = 14'd2013;
            {7'd61,7'd34}:		p = 14'd2074;
            {7'd61,7'd35}:		p = 14'd2135;
            {7'd61,7'd36}:		p = 14'd2196;
            {7'd61,7'd37}:		p = 14'd2257;
            {7'd61,7'd38}:		p = 14'd2318;
            {7'd61,7'd39}:		p = 14'd2379;
            {7'd61,7'd40}:		p = 14'd2440;
            {7'd61,7'd41}:		p = 14'd2501;
            {7'd61,7'd42}:		p = 14'd2562;
            {7'd61,7'd43}:		p = 14'd2623;
            {7'd61,7'd44}:		p = 14'd2684;
            {7'd61,7'd45}:		p = 14'd2745;
            {7'd61,7'd46}:		p = 14'd2806;
            {7'd61,7'd47}:		p = 14'd2867;
            {7'd61,7'd48}:		p = 14'd2928;
            {7'd61,7'd49}:		p = 14'd2989;
            {7'd61,7'd50}:		p = 14'd3050;
            {7'd61,7'd51}:		p = 14'd3111;
            {7'd61,7'd52}:		p = 14'd3172;
            {7'd61,7'd53}:		p = 14'd3233;
            {7'd61,7'd54}:		p = 14'd3294;
            {7'd61,7'd55}:		p = 14'd3355;
            {7'd61,7'd56}:		p = 14'd3416;
            {7'd61,7'd57}:		p = 14'd3477;
            {7'd61,7'd58}:		p = 14'd3538;
            {7'd61,7'd59}:		p = 14'd3599;
            {7'd61,7'd60}:		p = 14'd3660;
            {7'd61,7'd61}:		p = 14'd3721;
            {7'd61,7'd62}:		p = 14'd3782;
            {7'd61,7'd63}:		p = 14'd3843;
            {7'd61,7'd64}:		p = 14'd3904;
            {7'd61,7'd65}:		p = 14'd3965;
            {7'd61,7'd66}:		p = 14'd4026;
            {7'd61,7'd67}:		p = 14'd4087;
            {7'd61,7'd68}:		p = 14'd4148;
            {7'd61,7'd69}:		p = 14'd4209;
            {7'd61,7'd70}:		p = 14'd4270;
            {7'd61,7'd71}:		p = 14'd4331;
            {7'd61,7'd72}:		p = 14'd4392;
            {7'd61,7'd73}:		p = 14'd4453;
            {7'd61,7'd74}:		p = 14'd4514;
            {7'd61,7'd75}:		p = 14'd4575;
            {7'd61,7'd76}:		p = 14'd4636;
            {7'd61,7'd77}:		p = 14'd4697;
            {7'd61,7'd78}:		p = 14'd4758;
            {7'd61,7'd79}:		p = 14'd4819;
            {7'd61,7'd80}:		p = 14'd4880;
            {7'd61,7'd81}:		p = 14'd4941;
            {7'd61,7'd82}:		p = 14'd5002;
            {7'd61,7'd83}:		p = 14'd5063;
            {7'd61,7'd84}:		p = 14'd5124;
            {7'd61,7'd85}:		p = 14'd5185;
            {7'd61,7'd86}:		p = 14'd5246;
            {7'd61,7'd87}:		p = 14'd5307;
            {7'd61,7'd88}:		p = 14'd5368;
            {7'd61,7'd89}:		p = 14'd5429;
            {7'd61,7'd90}:		p = 14'd5490;
            {7'd61,7'd91}:		p = 14'd5551;
            {7'd61,7'd92}:		p = 14'd5612;
            {7'd61,7'd93}:		p = 14'd5673;
            {7'd61,7'd94}:		p = 14'd5734;
            {7'd61,7'd95}:		p = 14'd5795;
            {7'd61,7'd96}:		p = 14'd5856;
            {7'd61,7'd97}:		p = 14'd5917;
            {7'd61,7'd98}:		p = 14'd5978;
            {7'd61,7'd99}:		p = 14'd6039;
            {7'd61,7'd100}:		p = 14'd6100;
            {7'd61,7'd101}:		p = 14'd6161;
            {7'd61,7'd102}:		p = 14'd6222;
            {7'd61,7'd103}:		p = 14'd6283;
            {7'd61,7'd104}:		p = 14'd6344;
            {7'd61,7'd105}:		p = 14'd6405;
            {7'd61,7'd106}:		p = 14'd6466;
            {7'd61,7'd107}:		p = 14'd6527;
            {7'd61,7'd108}:		p = 14'd6588;
            {7'd61,7'd109}:		p = 14'd6649;
            {7'd61,7'd110}:		p = 14'd6710;
            {7'd61,7'd111}:		p = 14'd6771;
            {7'd61,7'd112}:		p = 14'd6832;
            {7'd61,7'd113}:		p = 14'd6893;
            {7'd61,7'd114}:		p = 14'd6954;
            {7'd61,7'd115}:		p = 14'd7015;
            {7'd61,7'd116}:		p = 14'd7076;
            {7'd61,7'd117}:		p = 14'd7137;
            {7'd61,7'd118}:		p = 14'd7198;
            {7'd61,7'd119}:		p = 14'd7259;
            {7'd61,7'd120}:		p = 14'd7320;
            {7'd61,7'd121}:		p = 14'd7381;
            {7'd61,7'd122}:		p = 14'd7442;
            {7'd61,7'd123}:		p = 14'd7503;
            {7'd61,7'd124}:		p = 14'd7564;
            {7'd61,7'd125}:		p = 14'd7625;
            {7'd61,7'd126}:		p = 14'd7686;
            {7'd61,7'd127}:		p = 14'd7747;
            {7'd62,7'd0}:		p = 14'd0;
            {7'd62,7'd1}:		p = 14'd62;
            {7'd62,7'd2}:		p = 14'd124;
            {7'd62,7'd3}:		p = 14'd186;
            {7'd62,7'd4}:		p = 14'd248;
            {7'd62,7'd5}:		p = 14'd310;
            {7'd62,7'd6}:		p = 14'd372;
            {7'd62,7'd7}:		p = 14'd434;
            {7'd62,7'd8}:		p = 14'd496;
            {7'd62,7'd9}:		p = 14'd558;
            {7'd62,7'd10}:		p = 14'd620;
            {7'd62,7'd11}:		p = 14'd682;
            {7'd62,7'd12}:		p = 14'd744;
            {7'd62,7'd13}:		p = 14'd806;
            {7'd62,7'd14}:		p = 14'd868;
            {7'd62,7'd15}:		p = 14'd930;
            {7'd62,7'd16}:		p = 14'd992;
            {7'd62,7'd17}:		p = 14'd1054;
            {7'd62,7'd18}:		p = 14'd1116;
            {7'd62,7'd19}:		p = 14'd1178;
            {7'd62,7'd20}:		p = 14'd1240;
            {7'd62,7'd21}:		p = 14'd1302;
            {7'd62,7'd22}:		p = 14'd1364;
            {7'd62,7'd23}:		p = 14'd1426;
            {7'd62,7'd24}:		p = 14'd1488;
            {7'd62,7'd25}:		p = 14'd1550;
            {7'd62,7'd26}:		p = 14'd1612;
            {7'd62,7'd27}:		p = 14'd1674;
            {7'd62,7'd28}:		p = 14'd1736;
            {7'd62,7'd29}:		p = 14'd1798;
            {7'd62,7'd30}:		p = 14'd1860;
            {7'd62,7'd31}:		p = 14'd1922;
            {7'd62,7'd32}:		p = 14'd1984;
            {7'd62,7'd33}:		p = 14'd2046;
            {7'd62,7'd34}:		p = 14'd2108;
            {7'd62,7'd35}:		p = 14'd2170;
            {7'd62,7'd36}:		p = 14'd2232;
            {7'd62,7'd37}:		p = 14'd2294;
            {7'd62,7'd38}:		p = 14'd2356;
            {7'd62,7'd39}:		p = 14'd2418;
            {7'd62,7'd40}:		p = 14'd2480;
            {7'd62,7'd41}:		p = 14'd2542;
            {7'd62,7'd42}:		p = 14'd2604;
            {7'd62,7'd43}:		p = 14'd2666;
            {7'd62,7'd44}:		p = 14'd2728;
            {7'd62,7'd45}:		p = 14'd2790;
            {7'd62,7'd46}:		p = 14'd2852;
            {7'd62,7'd47}:		p = 14'd2914;
            {7'd62,7'd48}:		p = 14'd2976;
            {7'd62,7'd49}:		p = 14'd3038;
            {7'd62,7'd50}:		p = 14'd3100;
            {7'd62,7'd51}:		p = 14'd3162;
            {7'd62,7'd52}:		p = 14'd3224;
            {7'd62,7'd53}:		p = 14'd3286;
            {7'd62,7'd54}:		p = 14'd3348;
            {7'd62,7'd55}:		p = 14'd3410;
            {7'd62,7'd56}:		p = 14'd3472;
            {7'd62,7'd57}:		p = 14'd3534;
            {7'd62,7'd58}:		p = 14'd3596;
            {7'd62,7'd59}:		p = 14'd3658;
            {7'd62,7'd60}:		p = 14'd3720;
            {7'd62,7'd61}:		p = 14'd3782;
            {7'd62,7'd62}:		p = 14'd3844;
            {7'd62,7'd63}:		p = 14'd3906;
            {7'd62,7'd64}:		p = 14'd3968;
            {7'd62,7'd65}:		p = 14'd4030;
            {7'd62,7'd66}:		p = 14'd4092;
            {7'd62,7'd67}:		p = 14'd4154;
            {7'd62,7'd68}:		p = 14'd4216;
            {7'd62,7'd69}:		p = 14'd4278;
            {7'd62,7'd70}:		p = 14'd4340;
            {7'd62,7'd71}:		p = 14'd4402;
            {7'd62,7'd72}:		p = 14'd4464;
            {7'd62,7'd73}:		p = 14'd4526;
            {7'd62,7'd74}:		p = 14'd4588;
            {7'd62,7'd75}:		p = 14'd4650;
            {7'd62,7'd76}:		p = 14'd4712;
            {7'd62,7'd77}:		p = 14'd4774;
            {7'd62,7'd78}:		p = 14'd4836;
            {7'd62,7'd79}:		p = 14'd4898;
            {7'd62,7'd80}:		p = 14'd4960;
            {7'd62,7'd81}:		p = 14'd5022;
            {7'd62,7'd82}:		p = 14'd5084;
            {7'd62,7'd83}:		p = 14'd5146;
            {7'd62,7'd84}:		p = 14'd5208;
            {7'd62,7'd85}:		p = 14'd5270;
            {7'd62,7'd86}:		p = 14'd5332;
            {7'd62,7'd87}:		p = 14'd5394;
            {7'd62,7'd88}:		p = 14'd5456;
            {7'd62,7'd89}:		p = 14'd5518;
            {7'd62,7'd90}:		p = 14'd5580;
            {7'd62,7'd91}:		p = 14'd5642;
            {7'd62,7'd92}:		p = 14'd5704;
            {7'd62,7'd93}:		p = 14'd5766;
            {7'd62,7'd94}:		p = 14'd5828;
            {7'd62,7'd95}:		p = 14'd5890;
            {7'd62,7'd96}:		p = 14'd5952;
            {7'd62,7'd97}:		p = 14'd6014;
            {7'd62,7'd98}:		p = 14'd6076;
            {7'd62,7'd99}:		p = 14'd6138;
            {7'd62,7'd100}:		p = 14'd6200;
            {7'd62,7'd101}:		p = 14'd6262;
            {7'd62,7'd102}:		p = 14'd6324;
            {7'd62,7'd103}:		p = 14'd6386;
            {7'd62,7'd104}:		p = 14'd6448;
            {7'd62,7'd105}:		p = 14'd6510;
            {7'd62,7'd106}:		p = 14'd6572;
            {7'd62,7'd107}:		p = 14'd6634;
            {7'd62,7'd108}:		p = 14'd6696;
            {7'd62,7'd109}:		p = 14'd6758;
            {7'd62,7'd110}:		p = 14'd6820;
            {7'd62,7'd111}:		p = 14'd6882;
            {7'd62,7'd112}:		p = 14'd6944;
            {7'd62,7'd113}:		p = 14'd7006;
            {7'd62,7'd114}:		p = 14'd7068;
            {7'd62,7'd115}:		p = 14'd7130;
            {7'd62,7'd116}:		p = 14'd7192;
            {7'd62,7'd117}:		p = 14'd7254;
            {7'd62,7'd118}:		p = 14'd7316;
            {7'd62,7'd119}:		p = 14'd7378;
            {7'd62,7'd120}:		p = 14'd7440;
            {7'd62,7'd121}:		p = 14'd7502;
            {7'd62,7'd122}:		p = 14'd7564;
            {7'd62,7'd123}:		p = 14'd7626;
            {7'd62,7'd124}:		p = 14'd7688;
            {7'd62,7'd125}:		p = 14'd7750;
            {7'd62,7'd126}:		p = 14'd7812;
            {7'd62,7'd127}:		p = 14'd7874;
            {7'd63,7'd0}:		p = 14'd0;
            {7'd63,7'd1}:		p = 14'd63;
            {7'd63,7'd2}:		p = 14'd126;
            {7'd63,7'd3}:		p = 14'd189;
            {7'd63,7'd4}:		p = 14'd252;
            {7'd63,7'd5}:		p = 14'd315;
            {7'd63,7'd6}:		p = 14'd378;
            {7'd63,7'd7}:		p = 14'd441;
            {7'd63,7'd8}:		p = 14'd504;
            {7'd63,7'd9}:		p = 14'd567;
            {7'd63,7'd10}:		p = 14'd630;
            {7'd63,7'd11}:		p = 14'd693;
            {7'd63,7'd12}:		p = 14'd756;
            {7'd63,7'd13}:		p = 14'd819;
            {7'd63,7'd14}:		p = 14'd882;
            {7'd63,7'd15}:		p = 14'd945;
            {7'd63,7'd16}:		p = 14'd1008;
            {7'd63,7'd17}:		p = 14'd1071;
            {7'd63,7'd18}:		p = 14'd1134;
            {7'd63,7'd19}:		p = 14'd1197;
            {7'd63,7'd20}:		p = 14'd1260;
            {7'd63,7'd21}:		p = 14'd1323;
            {7'd63,7'd22}:		p = 14'd1386;
            {7'd63,7'd23}:		p = 14'd1449;
            {7'd63,7'd24}:		p = 14'd1512;
            {7'd63,7'd25}:		p = 14'd1575;
            {7'd63,7'd26}:		p = 14'd1638;
            {7'd63,7'd27}:		p = 14'd1701;
            {7'd63,7'd28}:		p = 14'd1764;
            {7'd63,7'd29}:		p = 14'd1827;
            {7'd63,7'd30}:		p = 14'd1890;
            {7'd63,7'd31}:		p = 14'd1953;
            {7'd63,7'd32}:		p = 14'd2016;
            {7'd63,7'd33}:		p = 14'd2079;
            {7'd63,7'd34}:		p = 14'd2142;
            {7'd63,7'd35}:		p = 14'd2205;
            {7'd63,7'd36}:		p = 14'd2268;
            {7'd63,7'd37}:		p = 14'd2331;
            {7'd63,7'd38}:		p = 14'd2394;
            {7'd63,7'd39}:		p = 14'd2457;
            {7'd63,7'd40}:		p = 14'd2520;
            {7'd63,7'd41}:		p = 14'd2583;
            {7'd63,7'd42}:		p = 14'd2646;
            {7'd63,7'd43}:		p = 14'd2709;
            {7'd63,7'd44}:		p = 14'd2772;
            {7'd63,7'd45}:		p = 14'd2835;
            {7'd63,7'd46}:		p = 14'd2898;
            {7'd63,7'd47}:		p = 14'd2961;
            {7'd63,7'd48}:		p = 14'd3024;
            {7'd63,7'd49}:		p = 14'd3087;
            {7'd63,7'd50}:		p = 14'd3150;
            {7'd63,7'd51}:		p = 14'd3213;
            {7'd63,7'd52}:		p = 14'd3276;
            {7'd63,7'd53}:		p = 14'd3339;
            {7'd63,7'd54}:		p = 14'd3402;
            {7'd63,7'd55}:		p = 14'd3465;
            {7'd63,7'd56}:		p = 14'd3528;
            {7'd63,7'd57}:		p = 14'd3591;
            {7'd63,7'd58}:		p = 14'd3654;
            {7'd63,7'd59}:		p = 14'd3717;
            {7'd63,7'd60}:		p = 14'd3780;
            {7'd63,7'd61}:		p = 14'd3843;
            {7'd63,7'd62}:		p = 14'd3906;
            {7'd63,7'd63}:		p = 14'd3969;
            {7'd63,7'd64}:		p = 14'd4032;
            {7'd63,7'd65}:		p = 14'd4095;
            {7'd63,7'd66}:		p = 14'd4158;
            {7'd63,7'd67}:		p = 14'd4221;
            {7'd63,7'd68}:		p = 14'd4284;
            {7'd63,7'd69}:		p = 14'd4347;
            {7'd63,7'd70}:		p = 14'd4410;
            {7'd63,7'd71}:		p = 14'd4473;
            {7'd63,7'd72}:		p = 14'd4536;
            {7'd63,7'd73}:		p = 14'd4599;
            {7'd63,7'd74}:		p = 14'd4662;
            {7'd63,7'd75}:		p = 14'd4725;
            {7'd63,7'd76}:		p = 14'd4788;
            {7'd63,7'd77}:		p = 14'd4851;
            {7'd63,7'd78}:		p = 14'd4914;
            {7'd63,7'd79}:		p = 14'd4977;
            {7'd63,7'd80}:		p = 14'd5040;
            {7'd63,7'd81}:		p = 14'd5103;
            {7'd63,7'd82}:		p = 14'd5166;
            {7'd63,7'd83}:		p = 14'd5229;
            {7'd63,7'd84}:		p = 14'd5292;
            {7'd63,7'd85}:		p = 14'd5355;
            {7'd63,7'd86}:		p = 14'd5418;
            {7'd63,7'd87}:		p = 14'd5481;
            {7'd63,7'd88}:		p = 14'd5544;
            {7'd63,7'd89}:		p = 14'd5607;
            {7'd63,7'd90}:		p = 14'd5670;
            {7'd63,7'd91}:		p = 14'd5733;
            {7'd63,7'd92}:		p = 14'd5796;
            {7'd63,7'd93}:		p = 14'd5859;
            {7'd63,7'd94}:		p = 14'd5922;
            {7'd63,7'd95}:		p = 14'd5985;
            {7'd63,7'd96}:		p = 14'd6048;
            {7'd63,7'd97}:		p = 14'd6111;
            {7'd63,7'd98}:		p = 14'd6174;
            {7'd63,7'd99}:		p = 14'd6237;
            {7'd63,7'd100}:		p = 14'd6300;
            {7'd63,7'd101}:		p = 14'd6363;
            {7'd63,7'd102}:		p = 14'd6426;
            {7'd63,7'd103}:		p = 14'd6489;
            {7'd63,7'd104}:		p = 14'd6552;
            {7'd63,7'd105}:		p = 14'd6615;
            {7'd63,7'd106}:		p = 14'd6678;
            {7'd63,7'd107}:		p = 14'd6741;
            {7'd63,7'd108}:		p = 14'd6804;
            {7'd63,7'd109}:		p = 14'd6867;
            {7'd63,7'd110}:		p = 14'd6930;
            {7'd63,7'd111}:		p = 14'd6993;
            {7'd63,7'd112}:		p = 14'd7056;
            {7'd63,7'd113}:		p = 14'd7119;
            {7'd63,7'd114}:		p = 14'd7182;
            {7'd63,7'd115}:		p = 14'd7245;
            {7'd63,7'd116}:		p = 14'd7308;
            {7'd63,7'd117}:		p = 14'd7371;
            {7'd63,7'd118}:		p = 14'd7434;
            {7'd63,7'd119}:		p = 14'd7497;
            {7'd63,7'd120}:		p = 14'd7560;
            {7'd63,7'd121}:		p = 14'd7623;
            {7'd63,7'd122}:		p = 14'd7686;
            {7'd63,7'd123}:		p = 14'd7749;
            {7'd63,7'd124}:		p = 14'd7812;
            {7'd63,7'd125}:		p = 14'd7875;
            {7'd63,7'd126}:		p = 14'd7938;
            {7'd63,7'd127}:		p = 14'd8001;
            {7'd64,7'd0}:		p = 14'd0;
            {7'd64,7'd1}:		p = 14'd64;
            {7'd64,7'd2}:		p = 14'd128;
            {7'd64,7'd3}:		p = 14'd192;
            {7'd64,7'd4}:		p = 14'd256;
            {7'd64,7'd5}:		p = 14'd320;
            {7'd64,7'd6}:		p = 14'd384;
            {7'd64,7'd7}:		p = 14'd448;
            {7'd64,7'd8}:		p = 14'd512;
            {7'd64,7'd9}:		p = 14'd576;
            {7'd64,7'd10}:		p = 14'd640;
            {7'd64,7'd11}:		p = 14'd704;
            {7'd64,7'd12}:		p = 14'd768;
            {7'd64,7'd13}:		p = 14'd832;
            {7'd64,7'd14}:		p = 14'd896;
            {7'd64,7'd15}:		p = 14'd960;
            {7'd64,7'd16}:		p = 14'd1024;
            {7'd64,7'd17}:		p = 14'd1088;
            {7'd64,7'd18}:		p = 14'd1152;
            {7'd64,7'd19}:		p = 14'd1216;
            {7'd64,7'd20}:		p = 14'd1280;
            {7'd64,7'd21}:		p = 14'd1344;
            {7'd64,7'd22}:		p = 14'd1408;
            {7'd64,7'd23}:		p = 14'd1472;
            {7'd64,7'd24}:		p = 14'd1536;
            {7'd64,7'd25}:		p = 14'd1600;
            {7'd64,7'd26}:		p = 14'd1664;
            {7'd64,7'd27}:		p = 14'd1728;
            {7'd64,7'd28}:		p = 14'd1792;
            {7'd64,7'd29}:		p = 14'd1856;
            {7'd64,7'd30}:		p = 14'd1920;
            {7'd64,7'd31}:		p = 14'd1984;
            {7'd64,7'd32}:		p = 14'd2048;
            {7'd64,7'd33}:		p = 14'd2112;
            {7'd64,7'd34}:		p = 14'd2176;
            {7'd64,7'd35}:		p = 14'd2240;
            {7'd64,7'd36}:		p = 14'd2304;
            {7'd64,7'd37}:		p = 14'd2368;
            {7'd64,7'd38}:		p = 14'd2432;
            {7'd64,7'd39}:		p = 14'd2496;
            {7'd64,7'd40}:		p = 14'd2560;
            {7'd64,7'd41}:		p = 14'd2624;
            {7'd64,7'd42}:		p = 14'd2688;
            {7'd64,7'd43}:		p = 14'd2752;
            {7'd64,7'd44}:		p = 14'd2816;
            {7'd64,7'd45}:		p = 14'd2880;
            {7'd64,7'd46}:		p = 14'd2944;
            {7'd64,7'd47}:		p = 14'd3008;
            {7'd64,7'd48}:		p = 14'd3072;
            {7'd64,7'd49}:		p = 14'd3136;
            {7'd64,7'd50}:		p = 14'd3200;
            {7'd64,7'd51}:		p = 14'd3264;
            {7'd64,7'd52}:		p = 14'd3328;
            {7'd64,7'd53}:		p = 14'd3392;
            {7'd64,7'd54}:		p = 14'd3456;
            {7'd64,7'd55}:		p = 14'd3520;
            {7'd64,7'd56}:		p = 14'd3584;
            {7'd64,7'd57}:		p = 14'd3648;
            {7'd64,7'd58}:		p = 14'd3712;
            {7'd64,7'd59}:		p = 14'd3776;
            {7'd64,7'd60}:		p = 14'd3840;
            {7'd64,7'd61}:		p = 14'd3904;
            {7'd64,7'd62}:		p = 14'd3968;
            {7'd64,7'd63}:		p = 14'd4032;
            {7'd64,7'd64}:		p = 14'd4096;
            {7'd64,7'd65}:		p = 14'd4160;
            {7'd64,7'd66}:		p = 14'd4224;
            {7'd64,7'd67}:		p = 14'd4288;
            {7'd64,7'd68}:		p = 14'd4352;
            {7'd64,7'd69}:		p = 14'd4416;
            {7'd64,7'd70}:		p = 14'd4480;
            {7'd64,7'd71}:		p = 14'd4544;
            {7'd64,7'd72}:		p = 14'd4608;
            {7'd64,7'd73}:		p = 14'd4672;
            {7'd64,7'd74}:		p = 14'd4736;
            {7'd64,7'd75}:		p = 14'd4800;
            {7'd64,7'd76}:		p = 14'd4864;
            {7'd64,7'd77}:		p = 14'd4928;
            {7'd64,7'd78}:		p = 14'd4992;
            {7'd64,7'd79}:		p = 14'd5056;
            {7'd64,7'd80}:		p = 14'd5120;
            {7'd64,7'd81}:		p = 14'd5184;
            {7'd64,7'd82}:		p = 14'd5248;
            {7'd64,7'd83}:		p = 14'd5312;
            {7'd64,7'd84}:		p = 14'd5376;
            {7'd64,7'd85}:		p = 14'd5440;
            {7'd64,7'd86}:		p = 14'd5504;
            {7'd64,7'd87}:		p = 14'd5568;
            {7'd64,7'd88}:		p = 14'd5632;
            {7'd64,7'd89}:		p = 14'd5696;
            {7'd64,7'd90}:		p = 14'd5760;
            {7'd64,7'd91}:		p = 14'd5824;
            {7'd64,7'd92}:		p = 14'd5888;
            {7'd64,7'd93}:		p = 14'd5952;
            {7'd64,7'd94}:		p = 14'd6016;
            {7'd64,7'd95}:		p = 14'd6080;
            {7'd64,7'd96}:		p = 14'd6144;
            {7'd64,7'd97}:		p = 14'd6208;
            {7'd64,7'd98}:		p = 14'd6272;
            {7'd64,7'd99}:		p = 14'd6336;
            {7'd64,7'd100}:		p = 14'd6400;
            {7'd64,7'd101}:		p = 14'd6464;
            {7'd64,7'd102}:		p = 14'd6528;
            {7'd64,7'd103}:		p = 14'd6592;
            {7'd64,7'd104}:		p = 14'd6656;
            {7'd64,7'd105}:		p = 14'd6720;
            {7'd64,7'd106}:		p = 14'd6784;
            {7'd64,7'd107}:		p = 14'd6848;
            {7'd64,7'd108}:		p = 14'd6912;
            {7'd64,7'd109}:		p = 14'd6976;
            {7'd64,7'd110}:		p = 14'd7040;
            {7'd64,7'd111}:		p = 14'd7104;
            {7'd64,7'd112}:		p = 14'd7168;
            {7'd64,7'd113}:		p = 14'd7232;
            {7'd64,7'd114}:		p = 14'd7296;
            {7'd64,7'd115}:		p = 14'd7360;
            {7'd64,7'd116}:		p = 14'd7424;
            {7'd64,7'd117}:		p = 14'd7488;
            {7'd64,7'd118}:		p = 14'd7552;
            {7'd64,7'd119}:		p = 14'd7616;
            {7'd64,7'd120}:		p = 14'd7680;
            {7'd64,7'd121}:		p = 14'd7744;
            {7'd64,7'd122}:		p = 14'd7808;
            {7'd64,7'd123}:		p = 14'd7872;
            {7'd64,7'd124}:		p = 14'd7936;
            {7'd64,7'd125}:		p = 14'd8000;
            {7'd64,7'd126}:		p = 14'd8064;
            {7'd64,7'd127}:		p = 14'd8128;
            {7'd65,7'd0}:		p = 14'd0;
            {7'd65,7'd1}:		p = 14'd65;
            {7'd65,7'd2}:		p = 14'd130;
            {7'd65,7'd3}:		p = 14'd195;
            {7'd65,7'd4}:		p = 14'd260;
            {7'd65,7'd5}:		p = 14'd325;
            {7'd65,7'd6}:		p = 14'd390;
            {7'd65,7'd7}:		p = 14'd455;
            {7'd65,7'd8}:		p = 14'd520;
            {7'd65,7'd9}:		p = 14'd585;
            {7'd65,7'd10}:		p = 14'd650;
            {7'd65,7'd11}:		p = 14'd715;
            {7'd65,7'd12}:		p = 14'd780;
            {7'd65,7'd13}:		p = 14'd845;
            {7'd65,7'd14}:		p = 14'd910;
            {7'd65,7'd15}:		p = 14'd975;
            {7'd65,7'd16}:		p = 14'd1040;
            {7'd65,7'd17}:		p = 14'd1105;
            {7'd65,7'd18}:		p = 14'd1170;
            {7'd65,7'd19}:		p = 14'd1235;
            {7'd65,7'd20}:		p = 14'd1300;
            {7'd65,7'd21}:		p = 14'd1365;
            {7'd65,7'd22}:		p = 14'd1430;
            {7'd65,7'd23}:		p = 14'd1495;
            {7'd65,7'd24}:		p = 14'd1560;
            {7'd65,7'd25}:		p = 14'd1625;
            {7'd65,7'd26}:		p = 14'd1690;
            {7'd65,7'd27}:		p = 14'd1755;
            {7'd65,7'd28}:		p = 14'd1820;
            {7'd65,7'd29}:		p = 14'd1885;
            {7'd65,7'd30}:		p = 14'd1950;
            {7'd65,7'd31}:		p = 14'd2015;
            {7'd65,7'd32}:		p = 14'd2080;
            {7'd65,7'd33}:		p = 14'd2145;
            {7'd65,7'd34}:		p = 14'd2210;
            {7'd65,7'd35}:		p = 14'd2275;
            {7'd65,7'd36}:		p = 14'd2340;
            {7'd65,7'd37}:		p = 14'd2405;
            {7'd65,7'd38}:		p = 14'd2470;
            {7'd65,7'd39}:		p = 14'd2535;
            {7'd65,7'd40}:		p = 14'd2600;
            {7'd65,7'd41}:		p = 14'd2665;
            {7'd65,7'd42}:		p = 14'd2730;
            {7'd65,7'd43}:		p = 14'd2795;
            {7'd65,7'd44}:		p = 14'd2860;
            {7'd65,7'd45}:		p = 14'd2925;
            {7'd65,7'd46}:		p = 14'd2990;
            {7'd65,7'd47}:		p = 14'd3055;
            {7'd65,7'd48}:		p = 14'd3120;
            {7'd65,7'd49}:		p = 14'd3185;
            {7'd65,7'd50}:		p = 14'd3250;
            {7'd65,7'd51}:		p = 14'd3315;
            {7'd65,7'd52}:		p = 14'd3380;
            {7'd65,7'd53}:		p = 14'd3445;
            {7'd65,7'd54}:		p = 14'd3510;
            {7'd65,7'd55}:		p = 14'd3575;
            {7'd65,7'd56}:		p = 14'd3640;
            {7'd65,7'd57}:		p = 14'd3705;
            {7'd65,7'd58}:		p = 14'd3770;
            {7'd65,7'd59}:		p = 14'd3835;
            {7'd65,7'd60}:		p = 14'd3900;
            {7'd65,7'd61}:		p = 14'd3965;
            {7'd65,7'd62}:		p = 14'd4030;
            {7'd65,7'd63}:		p = 14'd4095;
            {7'd65,7'd64}:		p = 14'd4160;
            {7'd65,7'd65}:		p = 14'd4225;
            {7'd65,7'd66}:		p = 14'd4290;
            {7'd65,7'd67}:		p = 14'd4355;
            {7'd65,7'd68}:		p = 14'd4420;
            {7'd65,7'd69}:		p = 14'd4485;
            {7'd65,7'd70}:		p = 14'd4550;
            {7'd65,7'd71}:		p = 14'd4615;
            {7'd65,7'd72}:		p = 14'd4680;
            {7'd65,7'd73}:		p = 14'd4745;
            {7'd65,7'd74}:		p = 14'd4810;
            {7'd65,7'd75}:		p = 14'd4875;
            {7'd65,7'd76}:		p = 14'd4940;
            {7'd65,7'd77}:		p = 14'd5005;
            {7'd65,7'd78}:		p = 14'd5070;
            {7'd65,7'd79}:		p = 14'd5135;
            {7'd65,7'd80}:		p = 14'd5200;
            {7'd65,7'd81}:		p = 14'd5265;
            {7'd65,7'd82}:		p = 14'd5330;
            {7'd65,7'd83}:		p = 14'd5395;
            {7'd65,7'd84}:		p = 14'd5460;
            {7'd65,7'd85}:		p = 14'd5525;
            {7'd65,7'd86}:		p = 14'd5590;
            {7'd65,7'd87}:		p = 14'd5655;
            {7'd65,7'd88}:		p = 14'd5720;
            {7'd65,7'd89}:		p = 14'd5785;
            {7'd65,7'd90}:		p = 14'd5850;
            {7'd65,7'd91}:		p = 14'd5915;
            {7'd65,7'd92}:		p = 14'd5980;
            {7'd65,7'd93}:		p = 14'd6045;
            {7'd65,7'd94}:		p = 14'd6110;
            {7'd65,7'd95}:		p = 14'd6175;
            {7'd65,7'd96}:		p = 14'd6240;
            {7'd65,7'd97}:		p = 14'd6305;
            {7'd65,7'd98}:		p = 14'd6370;
            {7'd65,7'd99}:		p = 14'd6435;
            {7'd65,7'd100}:		p = 14'd6500;
            {7'd65,7'd101}:		p = 14'd6565;
            {7'd65,7'd102}:		p = 14'd6630;
            {7'd65,7'd103}:		p = 14'd6695;
            {7'd65,7'd104}:		p = 14'd6760;
            {7'd65,7'd105}:		p = 14'd6825;
            {7'd65,7'd106}:		p = 14'd6890;
            {7'd65,7'd107}:		p = 14'd6955;
            {7'd65,7'd108}:		p = 14'd7020;
            {7'd65,7'd109}:		p = 14'd7085;
            {7'd65,7'd110}:		p = 14'd7150;
            {7'd65,7'd111}:		p = 14'd7215;
            {7'd65,7'd112}:		p = 14'd7280;
            {7'd65,7'd113}:		p = 14'd7345;
            {7'd65,7'd114}:		p = 14'd7410;
            {7'd65,7'd115}:		p = 14'd7475;
            {7'd65,7'd116}:		p = 14'd7540;
            {7'd65,7'd117}:		p = 14'd7605;
            {7'd65,7'd118}:		p = 14'd7670;
            {7'd65,7'd119}:		p = 14'd7735;
            {7'd65,7'd120}:		p = 14'd7800;
            {7'd65,7'd121}:		p = 14'd7865;
            {7'd65,7'd122}:		p = 14'd7930;
            {7'd65,7'd123}:		p = 14'd7995;
            {7'd65,7'd124}:		p = 14'd8060;
            {7'd65,7'd125}:		p = 14'd8125;
            {7'd65,7'd126}:		p = 14'd8190;
            {7'd65,7'd127}:		p = 14'd8255;
            {7'd66,7'd0}:		p = 14'd0;
            {7'd66,7'd1}:		p = 14'd66;
            {7'd66,7'd2}:		p = 14'd132;
            {7'd66,7'd3}:		p = 14'd198;
            {7'd66,7'd4}:		p = 14'd264;
            {7'd66,7'd5}:		p = 14'd330;
            {7'd66,7'd6}:		p = 14'd396;
            {7'd66,7'd7}:		p = 14'd462;
            {7'd66,7'd8}:		p = 14'd528;
            {7'd66,7'd9}:		p = 14'd594;
            {7'd66,7'd10}:		p = 14'd660;
            {7'd66,7'd11}:		p = 14'd726;
            {7'd66,7'd12}:		p = 14'd792;
            {7'd66,7'd13}:		p = 14'd858;
            {7'd66,7'd14}:		p = 14'd924;
            {7'd66,7'd15}:		p = 14'd990;
            {7'd66,7'd16}:		p = 14'd1056;
            {7'd66,7'd17}:		p = 14'd1122;
            {7'd66,7'd18}:		p = 14'd1188;
            {7'd66,7'd19}:		p = 14'd1254;
            {7'd66,7'd20}:		p = 14'd1320;
            {7'd66,7'd21}:		p = 14'd1386;
            {7'd66,7'd22}:		p = 14'd1452;
            {7'd66,7'd23}:		p = 14'd1518;
            {7'd66,7'd24}:		p = 14'd1584;
            {7'd66,7'd25}:		p = 14'd1650;
            {7'd66,7'd26}:		p = 14'd1716;
            {7'd66,7'd27}:		p = 14'd1782;
            {7'd66,7'd28}:		p = 14'd1848;
            {7'd66,7'd29}:		p = 14'd1914;
            {7'd66,7'd30}:		p = 14'd1980;
            {7'd66,7'd31}:		p = 14'd2046;
            {7'd66,7'd32}:		p = 14'd2112;
            {7'd66,7'd33}:		p = 14'd2178;
            {7'd66,7'd34}:		p = 14'd2244;
            {7'd66,7'd35}:		p = 14'd2310;
            {7'd66,7'd36}:		p = 14'd2376;
            {7'd66,7'd37}:		p = 14'd2442;
            {7'd66,7'd38}:		p = 14'd2508;
            {7'd66,7'd39}:		p = 14'd2574;
            {7'd66,7'd40}:		p = 14'd2640;
            {7'd66,7'd41}:		p = 14'd2706;
            {7'd66,7'd42}:		p = 14'd2772;
            {7'd66,7'd43}:		p = 14'd2838;
            {7'd66,7'd44}:		p = 14'd2904;
            {7'd66,7'd45}:		p = 14'd2970;
            {7'd66,7'd46}:		p = 14'd3036;
            {7'd66,7'd47}:		p = 14'd3102;
            {7'd66,7'd48}:		p = 14'd3168;
            {7'd66,7'd49}:		p = 14'd3234;
            {7'd66,7'd50}:		p = 14'd3300;
            {7'd66,7'd51}:		p = 14'd3366;
            {7'd66,7'd52}:		p = 14'd3432;
            {7'd66,7'd53}:		p = 14'd3498;
            {7'd66,7'd54}:		p = 14'd3564;
            {7'd66,7'd55}:		p = 14'd3630;
            {7'd66,7'd56}:		p = 14'd3696;
            {7'd66,7'd57}:		p = 14'd3762;
            {7'd66,7'd58}:		p = 14'd3828;
            {7'd66,7'd59}:		p = 14'd3894;
            {7'd66,7'd60}:		p = 14'd3960;
            {7'd66,7'd61}:		p = 14'd4026;
            {7'd66,7'd62}:		p = 14'd4092;
            {7'd66,7'd63}:		p = 14'd4158;
            {7'd66,7'd64}:		p = 14'd4224;
            {7'd66,7'd65}:		p = 14'd4290;
            {7'd66,7'd66}:		p = 14'd4356;
            {7'd66,7'd67}:		p = 14'd4422;
            {7'd66,7'd68}:		p = 14'd4488;
            {7'd66,7'd69}:		p = 14'd4554;
            {7'd66,7'd70}:		p = 14'd4620;
            {7'd66,7'd71}:		p = 14'd4686;
            {7'd66,7'd72}:		p = 14'd4752;
            {7'd66,7'd73}:		p = 14'd4818;
            {7'd66,7'd74}:		p = 14'd4884;
            {7'd66,7'd75}:		p = 14'd4950;
            {7'd66,7'd76}:		p = 14'd5016;
            {7'd66,7'd77}:		p = 14'd5082;
            {7'd66,7'd78}:		p = 14'd5148;
            {7'd66,7'd79}:		p = 14'd5214;
            {7'd66,7'd80}:		p = 14'd5280;
            {7'd66,7'd81}:		p = 14'd5346;
            {7'd66,7'd82}:		p = 14'd5412;
            {7'd66,7'd83}:		p = 14'd5478;
            {7'd66,7'd84}:		p = 14'd5544;
            {7'd66,7'd85}:		p = 14'd5610;
            {7'd66,7'd86}:		p = 14'd5676;
            {7'd66,7'd87}:		p = 14'd5742;
            {7'd66,7'd88}:		p = 14'd5808;
            {7'd66,7'd89}:		p = 14'd5874;
            {7'd66,7'd90}:		p = 14'd5940;
            {7'd66,7'd91}:		p = 14'd6006;
            {7'd66,7'd92}:		p = 14'd6072;
            {7'd66,7'd93}:		p = 14'd6138;
            {7'd66,7'd94}:		p = 14'd6204;
            {7'd66,7'd95}:		p = 14'd6270;
            {7'd66,7'd96}:		p = 14'd6336;
            {7'd66,7'd97}:		p = 14'd6402;
            {7'd66,7'd98}:		p = 14'd6468;
            {7'd66,7'd99}:		p = 14'd6534;
            {7'd66,7'd100}:		p = 14'd6600;
            {7'd66,7'd101}:		p = 14'd6666;
            {7'd66,7'd102}:		p = 14'd6732;
            {7'd66,7'd103}:		p = 14'd6798;
            {7'd66,7'd104}:		p = 14'd6864;
            {7'd66,7'd105}:		p = 14'd6930;
            {7'd66,7'd106}:		p = 14'd6996;
            {7'd66,7'd107}:		p = 14'd7062;
            {7'd66,7'd108}:		p = 14'd7128;
            {7'd66,7'd109}:		p = 14'd7194;
            {7'd66,7'd110}:		p = 14'd7260;
            {7'd66,7'd111}:		p = 14'd7326;
            {7'd66,7'd112}:		p = 14'd7392;
            {7'd66,7'd113}:		p = 14'd7458;
            {7'd66,7'd114}:		p = 14'd7524;
            {7'd66,7'd115}:		p = 14'd7590;
            {7'd66,7'd116}:		p = 14'd7656;
            {7'd66,7'd117}:		p = 14'd7722;
            {7'd66,7'd118}:		p = 14'd7788;
            {7'd66,7'd119}:		p = 14'd7854;
            {7'd66,7'd120}:		p = 14'd7920;
            {7'd66,7'd121}:		p = 14'd7986;
            {7'd66,7'd122}:		p = 14'd8052;
            {7'd66,7'd123}:		p = 14'd8118;
            {7'd66,7'd124}:		p = 14'd8184;
            {7'd66,7'd125}:		p = 14'd8250;
            {7'd66,7'd126}:		p = 14'd8316;
            {7'd66,7'd127}:		p = 14'd8382;
            {7'd67,7'd0}:		p = 14'd0;
            {7'd67,7'd1}:		p = 14'd67;
            {7'd67,7'd2}:		p = 14'd134;
            {7'd67,7'd3}:		p = 14'd201;
            {7'd67,7'd4}:		p = 14'd268;
            {7'd67,7'd5}:		p = 14'd335;
            {7'd67,7'd6}:		p = 14'd402;
            {7'd67,7'd7}:		p = 14'd469;
            {7'd67,7'd8}:		p = 14'd536;
            {7'd67,7'd9}:		p = 14'd603;
            {7'd67,7'd10}:		p = 14'd670;
            {7'd67,7'd11}:		p = 14'd737;
            {7'd67,7'd12}:		p = 14'd804;
            {7'd67,7'd13}:		p = 14'd871;
            {7'd67,7'd14}:		p = 14'd938;
            {7'd67,7'd15}:		p = 14'd1005;
            {7'd67,7'd16}:		p = 14'd1072;
            {7'd67,7'd17}:		p = 14'd1139;
            {7'd67,7'd18}:		p = 14'd1206;
            {7'd67,7'd19}:		p = 14'd1273;
            {7'd67,7'd20}:		p = 14'd1340;
            {7'd67,7'd21}:		p = 14'd1407;
            {7'd67,7'd22}:		p = 14'd1474;
            {7'd67,7'd23}:		p = 14'd1541;
            {7'd67,7'd24}:		p = 14'd1608;
            {7'd67,7'd25}:		p = 14'd1675;
            {7'd67,7'd26}:		p = 14'd1742;
            {7'd67,7'd27}:		p = 14'd1809;
            {7'd67,7'd28}:		p = 14'd1876;
            {7'd67,7'd29}:		p = 14'd1943;
            {7'd67,7'd30}:		p = 14'd2010;
            {7'd67,7'd31}:		p = 14'd2077;
            {7'd67,7'd32}:		p = 14'd2144;
            {7'd67,7'd33}:		p = 14'd2211;
            {7'd67,7'd34}:		p = 14'd2278;
            {7'd67,7'd35}:		p = 14'd2345;
            {7'd67,7'd36}:		p = 14'd2412;
            {7'd67,7'd37}:		p = 14'd2479;
            {7'd67,7'd38}:		p = 14'd2546;
            {7'd67,7'd39}:		p = 14'd2613;
            {7'd67,7'd40}:		p = 14'd2680;
            {7'd67,7'd41}:		p = 14'd2747;
            {7'd67,7'd42}:		p = 14'd2814;
            {7'd67,7'd43}:		p = 14'd2881;
            {7'd67,7'd44}:		p = 14'd2948;
            {7'd67,7'd45}:		p = 14'd3015;
            {7'd67,7'd46}:		p = 14'd3082;
            {7'd67,7'd47}:		p = 14'd3149;
            {7'd67,7'd48}:		p = 14'd3216;
            {7'd67,7'd49}:		p = 14'd3283;
            {7'd67,7'd50}:		p = 14'd3350;
            {7'd67,7'd51}:		p = 14'd3417;
            {7'd67,7'd52}:		p = 14'd3484;
            {7'd67,7'd53}:		p = 14'd3551;
            {7'd67,7'd54}:		p = 14'd3618;
            {7'd67,7'd55}:		p = 14'd3685;
            {7'd67,7'd56}:		p = 14'd3752;
            {7'd67,7'd57}:		p = 14'd3819;
            {7'd67,7'd58}:		p = 14'd3886;
            {7'd67,7'd59}:		p = 14'd3953;
            {7'd67,7'd60}:		p = 14'd4020;
            {7'd67,7'd61}:		p = 14'd4087;
            {7'd67,7'd62}:		p = 14'd4154;
            {7'd67,7'd63}:		p = 14'd4221;
            {7'd67,7'd64}:		p = 14'd4288;
            {7'd67,7'd65}:		p = 14'd4355;
            {7'd67,7'd66}:		p = 14'd4422;
            {7'd67,7'd67}:		p = 14'd4489;
            {7'd67,7'd68}:		p = 14'd4556;
            {7'd67,7'd69}:		p = 14'd4623;
            {7'd67,7'd70}:		p = 14'd4690;
            {7'd67,7'd71}:		p = 14'd4757;
            {7'd67,7'd72}:		p = 14'd4824;
            {7'd67,7'd73}:		p = 14'd4891;
            {7'd67,7'd74}:		p = 14'd4958;
            {7'd67,7'd75}:		p = 14'd5025;
            {7'd67,7'd76}:		p = 14'd5092;
            {7'd67,7'd77}:		p = 14'd5159;
            {7'd67,7'd78}:		p = 14'd5226;
            {7'd67,7'd79}:		p = 14'd5293;
            {7'd67,7'd80}:		p = 14'd5360;
            {7'd67,7'd81}:		p = 14'd5427;
            {7'd67,7'd82}:		p = 14'd5494;
            {7'd67,7'd83}:		p = 14'd5561;
            {7'd67,7'd84}:		p = 14'd5628;
            {7'd67,7'd85}:		p = 14'd5695;
            {7'd67,7'd86}:		p = 14'd5762;
            {7'd67,7'd87}:		p = 14'd5829;
            {7'd67,7'd88}:		p = 14'd5896;
            {7'd67,7'd89}:		p = 14'd5963;
            {7'd67,7'd90}:		p = 14'd6030;
            {7'd67,7'd91}:		p = 14'd6097;
            {7'd67,7'd92}:		p = 14'd6164;
            {7'd67,7'd93}:		p = 14'd6231;
            {7'd67,7'd94}:		p = 14'd6298;
            {7'd67,7'd95}:		p = 14'd6365;
            {7'd67,7'd96}:		p = 14'd6432;
            {7'd67,7'd97}:		p = 14'd6499;
            {7'd67,7'd98}:		p = 14'd6566;
            {7'd67,7'd99}:		p = 14'd6633;
            {7'd67,7'd100}:		p = 14'd6700;
            {7'd67,7'd101}:		p = 14'd6767;
            {7'd67,7'd102}:		p = 14'd6834;
            {7'd67,7'd103}:		p = 14'd6901;
            {7'd67,7'd104}:		p = 14'd6968;
            {7'd67,7'd105}:		p = 14'd7035;
            {7'd67,7'd106}:		p = 14'd7102;
            {7'd67,7'd107}:		p = 14'd7169;
            {7'd67,7'd108}:		p = 14'd7236;
            {7'd67,7'd109}:		p = 14'd7303;
            {7'd67,7'd110}:		p = 14'd7370;
            {7'd67,7'd111}:		p = 14'd7437;
            {7'd67,7'd112}:		p = 14'd7504;
            {7'd67,7'd113}:		p = 14'd7571;
            {7'd67,7'd114}:		p = 14'd7638;
            {7'd67,7'd115}:		p = 14'd7705;
            {7'd67,7'd116}:		p = 14'd7772;
            {7'd67,7'd117}:		p = 14'd7839;
            {7'd67,7'd118}:		p = 14'd7906;
            {7'd67,7'd119}:		p = 14'd7973;
            {7'd67,7'd120}:		p = 14'd8040;
            {7'd67,7'd121}:		p = 14'd8107;
            {7'd67,7'd122}:		p = 14'd8174;
            {7'd67,7'd123}:		p = 14'd8241;
            {7'd67,7'd124}:		p = 14'd8308;
            {7'd67,7'd125}:		p = 14'd8375;
            {7'd67,7'd126}:		p = 14'd8442;
            {7'd67,7'd127}:		p = 14'd8509;
            {7'd68,7'd0}:		p = 14'd0;
            {7'd68,7'd1}:		p = 14'd68;
            {7'd68,7'd2}:		p = 14'd136;
            {7'd68,7'd3}:		p = 14'd204;
            {7'd68,7'd4}:		p = 14'd272;
            {7'd68,7'd5}:		p = 14'd340;
            {7'd68,7'd6}:		p = 14'd408;
            {7'd68,7'd7}:		p = 14'd476;
            {7'd68,7'd8}:		p = 14'd544;
            {7'd68,7'd9}:		p = 14'd612;
            {7'd68,7'd10}:		p = 14'd680;
            {7'd68,7'd11}:		p = 14'd748;
            {7'd68,7'd12}:		p = 14'd816;
            {7'd68,7'd13}:		p = 14'd884;
            {7'd68,7'd14}:		p = 14'd952;
            {7'd68,7'd15}:		p = 14'd1020;
            {7'd68,7'd16}:		p = 14'd1088;
            {7'd68,7'd17}:		p = 14'd1156;
            {7'd68,7'd18}:		p = 14'd1224;
            {7'd68,7'd19}:		p = 14'd1292;
            {7'd68,7'd20}:		p = 14'd1360;
            {7'd68,7'd21}:		p = 14'd1428;
            {7'd68,7'd22}:		p = 14'd1496;
            {7'd68,7'd23}:		p = 14'd1564;
            {7'd68,7'd24}:		p = 14'd1632;
            {7'd68,7'd25}:		p = 14'd1700;
            {7'd68,7'd26}:		p = 14'd1768;
            {7'd68,7'd27}:		p = 14'd1836;
            {7'd68,7'd28}:		p = 14'd1904;
            {7'd68,7'd29}:		p = 14'd1972;
            {7'd68,7'd30}:		p = 14'd2040;
            {7'd68,7'd31}:		p = 14'd2108;
            {7'd68,7'd32}:		p = 14'd2176;
            {7'd68,7'd33}:		p = 14'd2244;
            {7'd68,7'd34}:		p = 14'd2312;
            {7'd68,7'd35}:		p = 14'd2380;
            {7'd68,7'd36}:		p = 14'd2448;
            {7'd68,7'd37}:		p = 14'd2516;
            {7'd68,7'd38}:		p = 14'd2584;
            {7'd68,7'd39}:		p = 14'd2652;
            {7'd68,7'd40}:		p = 14'd2720;
            {7'd68,7'd41}:		p = 14'd2788;
            {7'd68,7'd42}:		p = 14'd2856;
            {7'd68,7'd43}:		p = 14'd2924;
            {7'd68,7'd44}:		p = 14'd2992;
            {7'd68,7'd45}:		p = 14'd3060;
            {7'd68,7'd46}:		p = 14'd3128;
            {7'd68,7'd47}:		p = 14'd3196;
            {7'd68,7'd48}:		p = 14'd3264;
            {7'd68,7'd49}:		p = 14'd3332;
            {7'd68,7'd50}:		p = 14'd3400;
            {7'd68,7'd51}:		p = 14'd3468;
            {7'd68,7'd52}:		p = 14'd3536;
            {7'd68,7'd53}:		p = 14'd3604;
            {7'd68,7'd54}:		p = 14'd3672;
            {7'd68,7'd55}:		p = 14'd3740;
            {7'd68,7'd56}:		p = 14'd3808;
            {7'd68,7'd57}:		p = 14'd3876;
            {7'd68,7'd58}:		p = 14'd3944;
            {7'd68,7'd59}:		p = 14'd4012;
            {7'd68,7'd60}:		p = 14'd4080;
            {7'd68,7'd61}:		p = 14'd4148;
            {7'd68,7'd62}:		p = 14'd4216;
            {7'd68,7'd63}:		p = 14'd4284;
            {7'd68,7'd64}:		p = 14'd4352;
            {7'd68,7'd65}:		p = 14'd4420;
            {7'd68,7'd66}:		p = 14'd4488;
            {7'd68,7'd67}:		p = 14'd4556;
            {7'd68,7'd68}:		p = 14'd4624;
            {7'd68,7'd69}:		p = 14'd4692;
            {7'd68,7'd70}:		p = 14'd4760;
            {7'd68,7'd71}:		p = 14'd4828;
            {7'd68,7'd72}:		p = 14'd4896;
            {7'd68,7'd73}:		p = 14'd4964;
            {7'd68,7'd74}:		p = 14'd5032;
            {7'd68,7'd75}:		p = 14'd5100;
            {7'd68,7'd76}:		p = 14'd5168;
            {7'd68,7'd77}:		p = 14'd5236;
            {7'd68,7'd78}:		p = 14'd5304;
            {7'd68,7'd79}:		p = 14'd5372;
            {7'd68,7'd80}:		p = 14'd5440;
            {7'd68,7'd81}:		p = 14'd5508;
            {7'd68,7'd82}:		p = 14'd5576;
            {7'd68,7'd83}:		p = 14'd5644;
            {7'd68,7'd84}:		p = 14'd5712;
            {7'd68,7'd85}:		p = 14'd5780;
            {7'd68,7'd86}:		p = 14'd5848;
            {7'd68,7'd87}:		p = 14'd5916;
            {7'd68,7'd88}:		p = 14'd5984;
            {7'd68,7'd89}:		p = 14'd6052;
            {7'd68,7'd90}:		p = 14'd6120;
            {7'd68,7'd91}:		p = 14'd6188;
            {7'd68,7'd92}:		p = 14'd6256;
            {7'd68,7'd93}:		p = 14'd6324;
            {7'd68,7'd94}:		p = 14'd6392;
            {7'd68,7'd95}:		p = 14'd6460;
            {7'd68,7'd96}:		p = 14'd6528;
            {7'd68,7'd97}:		p = 14'd6596;
            {7'd68,7'd98}:		p = 14'd6664;
            {7'd68,7'd99}:		p = 14'd6732;
            {7'd68,7'd100}:		p = 14'd6800;
            {7'd68,7'd101}:		p = 14'd6868;
            {7'd68,7'd102}:		p = 14'd6936;
            {7'd68,7'd103}:		p = 14'd7004;
            {7'd68,7'd104}:		p = 14'd7072;
            {7'd68,7'd105}:		p = 14'd7140;
            {7'd68,7'd106}:		p = 14'd7208;
            {7'd68,7'd107}:		p = 14'd7276;
            {7'd68,7'd108}:		p = 14'd7344;
            {7'd68,7'd109}:		p = 14'd7412;
            {7'd68,7'd110}:		p = 14'd7480;
            {7'd68,7'd111}:		p = 14'd7548;
            {7'd68,7'd112}:		p = 14'd7616;
            {7'd68,7'd113}:		p = 14'd7684;
            {7'd68,7'd114}:		p = 14'd7752;
            {7'd68,7'd115}:		p = 14'd7820;
            {7'd68,7'd116}:		p = 14'd7888;
            {7'd68,7'd117}:		p = 14'd7956;
            {7'd68,7'd118}:		p = 14'd8024;
            {7'd68,7'd119}:		p = 14'd8092;
            {7'd68,7'd120}:		p = 14'd8160;
            {7'd68,7'd121}:		p = 14'd8228;
            {7'd68,7'd122}:		p = 14'd8296;
            {7'd68,7'd123}:		p = 14'd8364;
            {7'd68,7'd124}:		p = 14'd8432;
            {7'd68,7'd125}:		p = 14'd8500;
            {7'd68,7'd126}:		p = 14'd8568;
            {7'd68,7'd127}:		p = 14'd8636;
            {7'd69,7'd0}:		p = 14'd0;
            {7'd69,7'd1}:		p = 14'd69;
            {7'd69,7'd2}:		p = 14'd138;
            {7'd69,7'd3}:		p = 14'd207;
            {7'd69,7'd4}:		p = 14'd276;
            {7'd69,7'd5}:		p = 14'd345;
            {7'd69,7'd6}:		p = 14'd414;
            {7'd69,7'd7}:		p = 14'd483;
            {7'd69,7'd8}:		p = 14'd552;
            {7'd69,7'd9}:		p = 14'd621;
            {7'd69,7'd10}:		p = 14'd690;
            {7'd69,7'd11}:		p = 14'd759;
            {7'd69,7'd12}:		p = 14'd828;
            {7'd69,7'd13}:		p = 14'd897;
            {7'd69,7'd14}:		p = 14'd966;
            {7'd69,7'd15}:		p = 14'd1035;
            {7'd69,7'd16}:		p = 14'd1104;
            {7'd69,7'd17}:		p = 14'd1173;
            {7'd69,7'd18}:		p = 14'd1242;
            {7'd69,7'd19}:		p = 14'd1311;
            {7'd69,7'd20}:		p = 14'd1380;
            {7'd69,7'd21}:		p = 14'd1449;
            {7'd69,7'd22}:		p = 14'd1518;
            {7'd69,7'd23}:		p = 14'd1587;
            {7'd69,7'd24}:		p = 14'd1656;
            {7'd69,7'd25}:		p = 14'd1725;
            {7'd69,7'd26}:		p = 14'd1794;
            {7'd69,7'd27}:		p = 14'd1863;
            {7'd69,7'd28}:		p = 14'd1932;
            {7'd69,7'd29}:		p = 14'd2001;
            {7'd69,7'd30}:		p = 14'd2070;
            {7'd69,7'd31}:		p = 14'd2139;
            {7'd69,7'd32}:		p = 14'd2208;
            {7'd69,7'd33}:		p = 14'd2277;
            {7'd69,7'd34}:		p = 14'd2346;
            {7'd69,7'd35}:		p = 14'd2415;
            {7'd69,7'd36}:		p = 14'd2484;
            {7'd69,7'd37}:		p = 14'd2553;
            {7'd69,7'd38}:		p = 14'd2622;
            {7'd69,7'd39}:		p = 14'd2691;
            {7'd69,7'd40}:		p = 14'd2760;
            {7'd69,7'd41}:		p = 14'd2829;
            {7'd69,7'd42}:		p = 14'd2898;
            {7'd69,7'd43}:		p = 14'd2967;
            {7'd69,7'd44}:		p = 14'd3036;
            {7'd69,7'd45}:		p = 14'd3105;
            {7'd69,7'd46}:		p = 14'd3174;
            {7'd69,7'd47}:		p = 14'd3243;
            {7'd69,7'd48}:		p = 14'd3312;
            {7'd69,7'd49}:		p = 14'd3381;
            {7'd69,7'd50}:		p = 14'd3450;
            {7'd69,7'd51}:		p = 14'd3519;
            {7'd69,7'd52}:		p = 14'd3588;
            {7'd69,7'd53}:		p = 14'd3657;
            {7'd69,7'd54}:		p = 14'd3726;
            {7'd69,7'd55}:		p = 14'd3795;
            {7'd69,7'd56}:		p = 14'd3864;
            {7'd69,7'd57}:		p = 14'd3933;
            {7'd69,7'd58}:		p = 14'd4002;
            {7'd69,7'd59}:		p = 14'd4071;
            {7'd69,7'd60}:		p = 14'd4140;
            {7'd69,7'd61}:		p = 14'd4209;
            {7'd69,7'd62}:		p = 14'd4278;
            {7'd69,7'd63}:		p = 14'd4347;
            {7'd69,7'd64}:		p = 14'd4416;
            {7'd69,7'd65}:		p = 14'd4485;
            {7'd69,7'd66}:		p = 14'd4554;
            {7'd69,7'd67}:		p = 14'd4623;
            {7'd69,7'd68}:		p = 14'd4692;
            {7'd69,7'd69}:		p = 14'd4761;
            {7'd69,7'd70}:		p = 14'd4830;
            {7'd69,7'd71}:		p = 14'd4899;
            {7'd69,7'd72}:		p = 14'd4968;
            {7'd69,7'd73}:		p = 14'd5037;
            {7'd69,7'd74}:		p = 14'd5106;
            {7'd69,7'd75}:		p = 14'd5175;
            {7'd69,7'd76}:		p = 14'd5244;
            {7'd69,7'd77}:		p = 14'd5313;
            {7'd69,7'd78}:		p = 14'd5382;
            {7'd69,7'd79}:		p = 14'd5451;
            {7'd69,7'd80}:		p = 14'd5520;
            {7'd69,7'd81}:		p = 14'd5589;
            {7'd69,7'd82}:		p = 14'd5658;
            {7'd69,7'd83}:		p = 14'd5727;
            {7'd69,7'd84}:		p = 14'd5796;
            {7'd69,7'd85}:		p = 14'd5865;
            {7'd69,7'd86}:		p = 14'd5934;
            {7'd69,7'd87}:		p = 14'd6003;
            {7'd69,7'd88}:		p = 14'd6072;
            {7'd69,7'd89}:		p = 14'd6141;
            {7'd69,7'd90}:		p = 14'd6210;
            {7'd69,7'd91}:		p = 14'd6279;
            {7'd69,7'd92}:		p = 14'd6348;
            {7'd69,7'd93}:		p = 14'd6417;
            {7'd69,7'd94}:		p = 14'd6486;
            {7'd69,7'd95}:		p = 14'd6555;
            {7'd69,7'd96}:		p = 14'd6624;
            {7'd69,7'd97}:		p = 14'd6693;
            {7'd69,7'd98}:		p = 14'd6762;
            {7'd69,7'd99}:		p = 14'd6831;
            {7'd69,7'd100}:		p = 14'd6900;
            {7'd69,7'd101}:		p = 14'd6969;
            {7'd69,7'd102}:		p = 14'd7038;
            {7'd69,7'd103}:		p = 14'd7107;
            {7'd69,7'd104}:		p = 14'd7176;
            {7'd69,7'd105}:		p = 14'd7245;
            {7'd69,7'd106}:		p = 14'd7314;
            {7'd69,7'd107}:		p = 14'd7383;
            {7'd69,7'd108}:		p = 14'd7452;
            {7'd69,7'd109}:		p = 14'd7521;
            {7'd69,7'd110}:		p = 14'd7590;
            {7'd69,7'd111}:		p = 14'd7659;
            {7'd69,7'd112}:		p = 14'd7728;
            {7'd69,7'd113}:		p = 14'd7797;
            {7'd69,7'd114}:		p = 14'd7866;
            {7'd69,7'd115}:		p = 14'd7935;
            {7'd69,7'd116}:		p = 14'd8004;
            {7'd69,7'd117}:		p = 14'd8073;
            {7'd69,7'd118}:		p = 14'd8142;
            {7'd69,7'd119}:		p = 14'd8211;
            {7'd69,7'd120}:		p = 14'd8280;
            {7'd69,7'd121}:		p = 14'd8349;
            {7'd69,7'd122}:		p = 14'd8418;
            {7'd69,7'd123}:		p = 14'd8487;
            {7'd69,7'd124}:		p = 14'd8556;
            {7'd69,7'd125}:		p = 14'd8625;
            {7'd69,7'd126}:		p = 14'd8694;
            {7'd69,7'd127}:		p = 14'd8763;
            {7'd70,7'd0}:		p = 14'd0;
            {7'd70,7'd1}:		p = 14'd70;
            {7'd70,7'd2}:		p = 14'd140;
            {7'd70,7'd3}:		p = 14'd210;
            {7'd70,7'd4}:		p = 14'd280;
            {7'd70,7'd5}:		p = 14'd350;
            {7'd70,7'd6}:		p = 14'd420;
            {7'd70,7'd7}:		p = 14'd490;
            {7'd70,7'd8}:		p = 14'd560;
            {7'd70,7'd9}:		p = 14'd630;
            {7'd70,7'd10}:		p = 14'd700;
            {7'd70,7'd11}:		p = 14'd770;
            {7'd70,7'd12}:		p = 14'd840;
            {7'd70,7'd13}:		p = 14'd910;
            {7'd70,7'd14}:		p = 14'd980;
            {7'd70,7'd15}:		p = 14'd1050;
            {7'd70,7'd16}:		p = 14'd1120;
            {7'd70,7'd17}:		p = 14'd1190;
            {7'd70,7'd18}:		p = 14'd1260;
            {7'd70,7'd19}:		p = 14'd1330;
            {7'd70,7'd20}:		p = 14'd1400;
            {7'd70,7'd21}:		p = 14'd1470;
            {7'd70,7'd22}:		p = 14'd1540;
            {7'd70,7'd23}:		p = 14'd1610;
            {7'd70,7'd24}:		p = 14'd1680;
            {7'd70,7'd25}:		p = 14'd1750;
            {7'd70,7'd26}:		p = 14'd1820;
            {7'd70,7'd27}:		p = 14'd1890;
            {7'd70,7'd28}:		p = 14'd1960;
            {7'd70,7'd29}:		p = 14'd2030;
            {7'd70,7'd30}:		p = 14'd2100;
            {7'd70,7'd31}:		p = 14'd2170;
            {7'd70,7'd32}:		p = 14'd2240;
            {7'd70,7'd33}:		p = 14'd2310;
            {7'd70,7'd34}:		p = 14'd2380;
            {7'd70,7'd35}:		p = 14'd2450;
            {7'd70,7'd36}:		p = 14'd2520;
            {7'd70,7'd37}:		p = 14'd2590;
            {7'd70,7'd38}:		p = 14'd2660;
            {7'd70,7'd39}:		p = 14'd2730;
            {7'd70,7'd40}:		p = 14'd2800;
            {7'd70,7'd41}:		p = 14'd2870;
            {7'd70,7'd42}:		p = 14'd2940;
            {7'd70,7'd43}:		p = 14'd3010;
            {7'd70,7'd44}:		p = 14'd3080;
            {7'd70,7'd45}:		p = 14'd3150;
            {7'd70,7'd46}:		p = 14'd3220;
            {7'd70,7'd47}:		p = 14'd3290;
            {7'd70,7'd48}:		p = 14'd3360;
            {7'd70,7'd49}:		p = 14'd3430;
            {7'd70,7'd50}:		p = 14'd3500;
            {7'd70,7'd51}:		p = 14'd3570;
            {7'd70,7'd52}:		p = 14'd3640;
            {7'd70,7'd53}:		p = 14'd3710;
            {7'd70,7'd54}:		p = 14'd3780;
            {7'd70,7'd55}:		p = 14'd3850;
            {7'd70,7'd56}:		p = 14'd3920;
            {7'd70,7'd57}:		p = 14'd3990;
            {7'd70,7'd58}:		p = 14'd4060;
            {7'd70,7'd59}:		p = 14'd4130;
            {7'd70,7'd60}:		p = 14'd4200;
            {7'd70,7'd61}:		p = 14'd4270;
            {7'd70,7'd62}:		p = 14'd4340;
            {7'd70,7'd63}:		p = 14'd4410;
            {7'd70,7'd64}:		p = 14'd4480;
            {7'd70,7'd65}:		p = 14'd4550;
            {7'd70,7'd66}:		p = 14'd4620;
            {7'd70,7'd67}:		p = 14'd4690;
            {7'd70,7'd68}:		p = 14'd4760;
            {7'd70,7'd69}:		p = 14'd4830;
            {7'd70,7'd70}:		p = 14'd4900;
            {7'd70,7'd71}:		p = 14'd4970;
            {7'd70,7'd72}:		p = 14'd5040;
            {7'd70,7'd73}:		p = 14'd5110;
            {7'd70,7'd74}:		p = 14'd5180;
            {7'd70,7'd75}:		p = 14'd5250;
            {7'd70,7'd76}:		p = 14'd5320;
            {7'd70,7'd77}:		p = 14'd5390;
            {7'd70,7'd78}:		p = 14'd5460;
            {7'd70,7'd79}:		p = 14'd5530;
            {7'd70,7'd80}:		p = 14'd5600;
            {7'd70,7'd81}:		p = 14'd5670;
            {7'd70,7'd82}:		p = 14'd5740;
            {7'd70,7'd83}:		p = 14'd5810;
            {7'd70,7'd84}:		p = 14'd5880;
            {7'd70,7'd85}:		p = 14'd5950;
            {7'd70,7'd86}:		p = 14'd6020;
            {7'd70,7'd87}:		p = 14'd6090;
            {7'd70,7'd88}:		p = 14'd6160;
            {7'd70,7'd89}:		p = 14'd6230;
            {7'd70,7'd90}:		p = 14'd6300;
            {7'd70,7'd91}:		p = 14'd6370;
            {7'd70,7'd92}:		p = 14'd6440;
            {7'd70,7'd93}:		p = 14'd6510;
            {7'd70,7'd94}:		p = 14'd6580;
            {7'd70,7'd95}:		p = 14'd6650;
            {7'd70,7'd96}:		p = 14'd6720;
            {7'd70,7'd97}:		p = 14'd6790;
            {7'd70,7'd98}:		p = 14'd6860;
            {7'd70,7'd99}:		p = 14'd6930;
            {7'd70,7'd100}:		p = 14'd7000;
            {7'd70,7'd101}:		p = 14'd7070;
            {7'd70,7'd102}:		p = 14'd7140;
            {7'd70,7'd103}:		p = 14'd7210;
            {7'd70,7'd104}:		p = 14'd7280;
            {7'd70,7'd105}:		p = 14'd7350;
            {7'd70,7'd106}:		p = 14'd7420;
            {7'd70,7'd107}:		p = 14'd7490;
            {7'd70,7'd108}:		p = 14'd7560;
            {7'd70,7'd109}:		p = 14'd7630;
            {7'd70,7'd110}:		p = 14'd7700;
            {7'd70,7'd111}:		p = 14'd7770;
            {7'd70,7'd112}:		p = 14'd7840;
            {7'd70,7'd113}:		p = 14'd7910;
            {7'd70,7'd114}:		p = 14'd7980;
            {7'd70,7'd115}:		p = 14'd8050;
            {7'd70,7'd116}:		p = 14'd8120;
            {7'd70,7'd117}:		p = 14'd8190;
            {7'd70,7'd118}:		p = 14'd8260;
            {7'd70,7'd119}:		p = 14'd8330;
            {7'd70,7'd120}:		p = 14'd8400;
            {7'd70,7'd121}:		p = 14'd8470;
            {7'd70,7'd122}:		p = 14'd8540;
            {7'd70,7'd123}:		p = 14'd8610;
            {7'd70,7'd124}:		p = 14'd8680;
            {7'd70,7'd125}:		p = 14'd8750;
            {7'd70,7'd126}:		p = 14'd8820;
            {7'd70,7'd127}:		p = 14'd8890;
            {7'd71,7'd0}:		p = 14'd0;
            {7'd71,7'd1}:		p = 14'd71;
            {7'd71,7'd2}:		p = 14'd142;
            {7'd71,7'd3}:		p = 14'd213;
            {7'd71,7'd4}:		p = 14'd284;
            {7'd71,7'd5}:		p = 14'd355;
            {7'd71,7'd6}:		p = 14'd426;
            {7'd71,7'd7}:		p = 14'd497;
            {7'd71,7'd8}:		p = 14'd568;
            {7'd71,7'd9}:		p = 14'd639;
            {7'd71,7'd10}:		p = 14'd710;
            {7'd71,7'd11}:		p = 14'd781;
            {7'd71,7'd12}:		p = 14'd852;
            {7'd71,7'd13}:		p = 14'd923;
            {7'd71,7'd14}:		p = 14'd994;
            {7'd71,7'd15}:		p = 14'd1065;
            {7'd71,7'd16}:		p = 14'd1136;
            {7'd71,7'd17}:		p = 14'd1207;
            {7'd71,7'd18}:		p = 14'd1278;
            {7'd71,7'd19}:		p = 14'd1349;
            {7'd71,7'd20}:		p = 14'd1420;
            {7'd71,7'd21}:		p = 14'd1491;
            {7'd71,7'd22}:		p = 14'd1562;
            {7'd71,7'd23}:		p = 14'd1633;
            {7'd71,7'd24}:		p = 14'd1704;
            {7'd71,7'd25}:		p = 14'd1775;
            {7'd71,7'd26}:		p = 14'd1846;
            {7'd71,7'd27}:		p = 14'd1917;
            {7'd71,7'd28}:		p = 14'd1988;
            {7'd71,7'd29}:		p = 14'd2059;
            {7'd71,7'd30}:		p = 14'd2130;
            {7'd71,7'd31}:		p = 14'd2201;
            {7'd71,7'd32}:		p = 14'd2272;
            {7'd71,7'd33}:		p = 14'd2343;
            {7'd71,7'd34}:		p = 14'd2414;
            {7'd71,7'd35}:		p = 14'd2485;
            {7'd71,7'd36}:		p = 14'd2556;
            {7'd71,7'd37}:		p = 14'd2627;
            {7'd71,7'd38}:		p = 14'd2698;
            {7'd71,7'd39}:		p = 14'd2769;
            {7'd71,7'd40}:		p = 14'd2840;
            {7'd71,7'd41}:		p = 14'd2911;
            {7'd71,7'd42}:		p = 14'd2982;
            {7'd71,7'd43}:		p = 14'd3053;
            {7'd71,7'd44}:		p = 14'd3124;
            {7'd71,7'd45}:		p = 14'd3195;
            {7'd71,7'd46}:		p = 14'd3266;
            {7'd71,7'd47}:		p = 14'd3337;
            {7'd71,7'd48}:		p = 14'd3408;
            {7'd71,7'd49}:		p = 14'd3479;
            {7'd71,7'd50}:		p = 14'd3550;
            {7'd71,7'd51}:		p = 14'd3621;
            {7'd71,7'd52}:		p = 14'd3692;
            {7'd71,7'd53}:		p = 14'd3763;
            {7'd71,7'd54}:		p = 14'd3834;
            {7'd71,7'd55}:		p = 14'd3905;
            {7'd71,7'd56}:		p = 14'd3976;
            {7'd71,7'd57}:		p = 14'd4047;
            {7'd71,7'd58}:		p = 14'd4118;
            {7'd71,7'd59}:		p = 14'd4189;
            {7'd71,7'd60}:		p = 14'd4260;
            {7'd71,7'd61}:		p = 14'd4331;
            {7'd71,7'd62}:		p = 14'd4402;
            {7'd71,7'd63}:		p = 14'd4473;
            {7'd71,7'd64}:		p = 14'd4544;
            {7'd71,7'd65}:		p = 14'd4615;
            {7'd71,7'd66}:		p = 14'd4686;
            {7'd71,7'd67}:		p = 14'd4757;
            {7'd71,7'd68}:		p = 14'd4828;
            {7'd71,7'd69}:		p = 14'd4899;
            {7'd71,7'd70}:		p = 14'd4970;
            {7'd71,7'd71}:		p = 14'd5041;
            {7'd71,7'd72}:		p = 14'd5112;
            {7'd71,7'd73}:		p = 14'd5183;
            {7'd71,7'd74}:		p = 14'd5254;
            {7'd71,7'd75}:		p = 14'd5325;
            {7'd71,7'd76}:		p = 14'd5396;
            {7'd71,7'd77}:		p = 14'd5467;
            {7'd71,7'd78}:		p = 14'd5538;
            {7'd71,7'd79}:		p = 14'd5609;
            {7'd71,7'd80}:		p = 14'd5680;
            {7'd71,7'd81}:		p = 14'd5751;
            {7'd71,7'd82}:		p = 14'd5822;
            {7'd71,7'd83}:		p = 14'd5893;
            {7'd71,7'd84}:		p = 14'd5964;
            {7'd71,7'd85}:		p = 14'd6035;
            {7'd71,7'd86}:		p = 14'd6106;
            {7'd71,7'd87}:		p = 14'd6177;
            {7'd71,7'd88}:		p = 14'd6248;
            {7'd71,7'd89}:		p = 14'd6319;
            {7'd71,7'd90}:		p = 14'd6390;
            {7'd71,7'd91}:		p = 14'd6461;
            {7'd71,7'd92}:		p = 14'd6532;
            {7'd71,7'd93}:		p = 14'd6603;
            {7'd71,7'd94}:		p = 14'd6674;
            {7'd71,7'd95}:		p = 14'd6745;
            {7'd71,7'd96}:		p = 14'd6816;
            {7'd71,7'd97}:		p = 14'd6887;
            {7'd71,7'd98}:		p = 14'd6958;
            {7'd71,7'd99}:		p = 14'd7029;
            {7'd71,7'd100}:		p = 14'd7100;
            {7'd71,7'd101}:		p = 14'd7171;
            {7'd71,7'd102}:		p = 14'd7242;
            {7'd71,7'd103}:		p = 14'd7313;
            {7'd71,7'd104}:		p = 14'd7384;
            {7'd71,7'd105}:		p = 14'd7455;
            {7'd71,7'd106}:		p = 14'd7526;
            {7'd71,7'd107}:		p = 14'd7597;
            {7'd71,7'd108}:		p = 14'd7668;
            {7'd71,7'd109}:		p = 14'd7739;
            {7'd71,7'd110}:		p = 14'd7810;
            {7'd71,7'd111}:		p = 14'd7881;
            {7'd71,7'd112}:		p = 14'd7952;
            {7'd71,7'd113}:		p = 14'd8023;
            {7'd71,7'd114}:		p = 14'd8094;
            {7'd71,7'd115}:		p = 14'd8165;
            {7'd71,7'd116}:		p = 14'd8236;
            {7'd71,7'd117}:		p = 14'd8307;
            {7'd71,7'd118}:		p = 14'd8378;
            {7'd71,7'd119}:		p = 14'd8449;
            {7'd71,7'd120}:		p = 14'd8520;
            {7'd71,7'd121}:		p = 14'd8591;
            {7'd71,7'd122}:		p = 14'd8662;
            {7'd71,7'd123}:		p = 14'd8733;
            {7'd71,7'd124}:		p = 14'd8804;
            {7'd71,7'd125}:		p = 14'd8875;
            {7'd71,7'd126}:		p = 14'd8946;
            {7'd71,7'd127}:		p = 14'd9017;
            {7'd72,7'd0}:		p = 14'd0;
            {7'd72,7'd1}:		p = 14'd72;
            {7'd72,7'd2}:		p = 14'd144;
            {7'd72,7'd3}:		p = 14'd216;
            {7'd72,7'd4}:		p = 14'd288;
            {7'd72,7'd5}:		p = 14'd360;
            {7'd72,7'd6}:		p = 14'd432;
            {7'd72,7'd7}:		p = 14'd504;
            {7'd72,7'd8}:		p = 14'd576;
            {7'd72,7'd9}:		p = 14'd648;
            {7'd72,7'd10}:		p = 14'd720;
            {7'd72,7'd11}:		p = 14'd792;
            {7'd72,7'd12}:		p = 14'd864;
            {7'd72,7'd13}:		p = 14'd936;
            {7'd72,7'd14}:		p = 14'd1008;
            {7'd72,7'd15}:		p = 14'd1080;
            {7'd72,7'd16}:		p = 14'd1152;
            {7'd72,7'd17}:		p = 14'd1224;
            {7'd72,7'd18}:		p = 14'd1296;
            {7'd72,7'd19}:		p = 14'd1368;
            {7'd72,7'd20}:		p = 14'd1440;
            {7'd72,7'd21}:		p = 14'd1512;
            {7'd72,7'd22}:		p = 14'd1584;
            {7'd72,7'd23}:		p = 14'd1656;
            {7'd72,7'd24}:		p = 14'd1728;
            {7'd72,7'd25}:		p = 14'd1800;
            {7'd72,7'd26}:		p = 14'd1872;
            {7'd72,7'd27}:		p = 14'd1944;
            {7'd72,7'd28}:		p = 14'd2016;
            {7'd72,7'd29}:		p = 14'd2088;
            {7'd72,7'd30}:		p = 14'd2160;
            {7'd72,7'd31}:		p = 14'd2232;
            {7'd72,7'd32}:		p = 14'd2304;
            {7'd72,7'd33}:		p = 14'd2376;
            {7'd72,7'd34}:		p = 14'd2448;
            {7'd72,7'd35}:		p = 14'd2520;
            {7'd72,7'd36}:		p = 14'd2592;
            {7'd72,7'd37}:		p = 14'd2664;
            {7'd72,7'd38}:		p = 14'd2736;
            {7'd72,7'd39}:		p = 14'd2808;
            {7'd72,7'd40}:		p = 14'd2880;
            {7'd72,7'd41}:		p = 14'd2952;
            {7'd72,7'd42}:		p = 14'd3024;
            {7'd72,7'd43}:		p = 14'd3096;
            {7'd72,7'd44}:		p = 14'd3168;
            {7'd72,7'd45}:		p = 14'd3240;
            {7'd72,7'd46}:		p = 14'd3312;
            {7'd72,7'd47}:		p = 14'd3384;
            {7'd72,7'd48}:		p = 14'd3456;
            {7'd72,7'd49}:		p = 14'd3528;
            {7'd72,7'd50}:		p = 14'd3600;
            {7'd72,7'd51}:		p = 14'd3672;
            {7'd72,7'd52}:		p = 14'd3744;
            {7'd72,7'd53}:		p = 14'd3816;
            {7'd72,7'd54}:		p = 14'd3888;
            {7'd72,7'd55}:		p = 14'd3960;
            {7'd72,7'd56}:		p = 14'd4032;
            {7'd72,7'd57}:		p = 14'd4104;
            {7'd72,7'd58}:		p = 14'd4176;
            {7'd72,7'd59}:		p = 14'd4248;
            {7'd72,7'd60}:		p = 14'd4320;
            {7'd72,7'd61}:		p = 14'd4392;
            {7'd72,7'd62}:		p = 14'd4464;
            {7'd72,7'd63}:		p = 14'd4536;
            {7'd72,7'd64}:		p = 14'd4608;
            {7'd72,7'd65}:		p = 14'd4680;
            {7'd72,7'd66}:		p = 14'd4752;
            {7'd72,7'd67}:		p = 14'd4824;
            {7'd72,7'd68}:		p = 14'd4896;
            {7'd72,7'd69}:		p = 14'd4968;
            {7'd72,7'd70}:		p = 14'd5040;
            {7'd72,7'd71}:		p = 14'd5112;
            {7'd72,7'd72}:		p = 14'd5184;
            {7'd72,7'd73}:		p = 14'd5256;
            {7'd72,7'd74}:		p = 14'd5328;
            {7'd72,7'd75}:		p = 14'd5400;
            {7'd72,7'd76}:		p = 14'd5472;
            {7'd72,7'd77}:		p = 14'd5544;
            {7'd72,7'd78}:		p = 14'd5616;
            {7'd72,7'd79}:		p = 14'd5688;
            {7'd72,7'd80}:		p = 14'd5760;
            {7'd72,7'd81}:		p = 14'd5832;
            {7'd72,7'd82}:		p = 14'd5904;
            {7'd72,7'd83}:		p = 14'd5976;
            {7'd72,7'd84}:		p = 14'd6048;
            {7'd72,7'd85}:		p = 14'd6120;
            {7'd72,7'd86}:		p = 14'd6192;
            {7'd72,7'd87}:		p = 14'd6264;
            {7'd72,7'd88}:		p = 14'd6336;
            {7'd72,7'd89}:		p = 14'd6408;
            {7'd72,7'd90}:		p = 14'd6480;
            {7'd72,7'd91}:		p = 14'd6552;
            {7'd72,7'd92}:		p = 14'd6624;
            {7'd72,7'd93}:		p = 14'd6696;
            {7'd72,7'd94}:		p = 14'd6768;
            {7'd72,7'd95}:		p = 14'd6840;
            {7'd72,7'd96}:		p = 14'd6912;
            {7'd72,7'd97}:		p = 14'd6984;
            {7'd72,7'd98}:		p = 14'd7056;
            {7'd72,7'd99}:		p = 14'd7128;
            {7'd72,7'd100}:		p = 14'd7200;
            {7'd72,7'd101}:		p = 14'd7272;
            {7'd72,7'd102}:		p = 14'd7344;
            {7'd72,7'd103}:		p = 14'd7416;
            {7'd72,7'd104}:		p = 14'd7488;
            {7'd72,7'd105}:		p = 14'd7560;
            {7'd72,7'd106}:		p = 14'd7632;
            {7'd72,7'd107}:		p = 14'd7704;
            {7'd72,7'd108}:		p = 14'd7776;
            {7'd72,7'd109}:		p = 14'd7848;
            {7'd72,7'd110}:		p = 14'd7920;
            {7'd72,7'd111}:		p = 14'd7992;
            {7'd72,7'd112}:		p = 14'd8064;
            {7'd72,7'd113}:		p = 14'd8136;
            {7'd72,7'd114}:		p = 14'd8208;
            {7'd72,7'd115}:		p = 14'd8280;
            {7'd72,7'd116}:		p = 14'd8352;
            {7'd72,7'd117}:		p = 14'd8424;
            {7'd72,7'd118}:		p = 14'd8496;
            {7'd72,7'd119}:		p = 14'd8568;
            {7'd72,7'd120}:		p = 14'd8640;
            {7'd72,7'd121}:		p = 14'd8712;
            {7'd72,7'd122}:		p = 14'd8784;
            {7'd72,7'd123}:		p = 14'd8856;
            {7'd72,7'd124}:		p = 14'd8928;
            {7'd72,7'd125}:		p = 14'd9000;
            {7'd72,7'd126}:		p = 14'd9072;
            {7'd72,7'd127}:		p = 14'd9144;
            {7'd73,7'd0}:		p = 14'd0;
            {7'd73,7'd1}:		p = 14'd73;
            {7'd73,7'd2}:		p = 14'd146;
            {7'd73,7'd3}:		p = 14'd219;
            {7'd73,7'd4}:		p = 14'd292;
            {7'd73,7'd5}:		p = 14'd365;
            {7'd73,7'd6}:		p = 14'd438;
            {7'd73,7'd7}:		p = 14'd511;
            {7'd73,7'd8}:		p = 14'd584;
            {7'd73,7'd9}:		p = 14'd657;
            {7'd73,7'd10}:		p = 14'd730;
            {7'd73,7'd11}:		p = 14'd803;
            {7'd73,7'd12}:		p = 14'd876;
            {7'd73,7'd13}:		p = 14'd949;
            {7'd73,7'd14}:		p = 14'd1022;
            {7'd73,7'd15}:		p = 14'd1095;
            {7'd73,7'd16}:		p = 14'd1168;
            {7'd73,7'd17}:		p = 14'd1241;
            {7'd73,7'd18}:		p = 14'd1314;
            {7'd73,7'd19}:		p = 14'd1387;
            {7'd73,7'd20}:		p = 14'd1460;
            {7'd73,7'd21}:		p = 14'd1533;
            {7'd73,7'd22}:		p = 14'd1606;
            {7'd73,7'd23}:		p = 14'd1679;
            {7'd73,7'd24}:		p = 14'd1752;
            {7'd73,7'd25}:		p = 14'd1825;
            {7'd73,7'd26}:		p = 14'd1898;
            {7'd73,7'd27}:		p = 14'd1971;
            {7'd73,7'd28}:		p = 14'd2044;
            {7'd73,7'd29}:		p = 14'd2117;
            {7'd73,7'd30}:		p = 14'd2190;
            {7'd73,7'd31}:		p = 14'd2263;
            {7'd73,7'd32}:		p = 14'd2336;
            {7'd73,7'd33}:		p = 14'd2409;
            {7'd73,7'd34}:		p = 14'd2482;
            {7'd73,7'd35}:		p = 14'd2555;
            {7'd73,7'd36}:		p = 14'd2628;
            {7'd73,7'd37}:		p = 14'd2701;
            {7'd73,7'd38}:		p = 14'd2774;
            {7'd73,7'd39}:		p = 14'd2847;
            {7'd73,7'd40}:		p = 14'd2920;
            {7'd73,7'd41}:		p = 14'd2993;
            {7'd73,7'd42}:		p = 14'd3066;
            {7'd73,7'd43}:		p = 14'd3139;
            {7'd73,7'd44}:		p = 14'd3212;
            {7'd73,7'd45}:		p = 14'd3285;
            {7'd73,7'd46}:		p = 14'd3358;
            {7'd73,7'd47}:		p = 14'd3431;
            {7'd73,7'd48}:		p = 14'd3504;
            {7'd73,7'd49}:		p = 14'd3577;
            {7'd73,7'd50}:		p = 14'd3650;
            {7'd73,7'd51}:		p = 14'd3723;
            {7'd73,7'd52}:		p = 14'd3796;
            {7'd73,7'd53}:		p = 14'd3869;
            {7'd73,7'd54}:		p = 14'd3942;
            {7'd73,7'd55}:		p = 14'd4015;
            {7'd73,7'd56}:		p = 14'd4088;
            {7'd73,7'd57}:		p = 14'd4161;
            {7'd73,7'd58}:		p = 14'd4234;
            {7'd73,7'd59}:		p = 14'd4307;
            {7'd73,7'd60}:		p = 14'd4380;
            {7'd73,7'd61}:		p = 14'd4453;
            {7'd73,7'd62}:		p = 14'd4526;
            {7'd73,7'd63}:		p = 14'd4599;
            {7'd73,7'd64}:		p = 14'd4672;
            {7'd73,7'd65}:		p = 14'd4745;
            {7'd73,7'd66}:		p = 14'd4818;
            {7'd73,7'd67}:		p = 14'd4891;
            {7'd73,7'd68}:		p = 14'd4964;
            {7'd73,7'd69}:		p = 14'd5037;
            {7'd73,7'd70}:		p = 14'd5110;
            {7'd73,7'd71}:		p = 14'd5183;
            {7'd73,7'd72}:		p = 14'd5256;
            {7'd73,7'd73}:		p = 14'd5329;
            {7'd73,7'd74}:		p = 14'd5402;
            {7'd73,7'd75}:		p = 14'd5475;
            {7'd73,7'd76}:		p = 14'd5548;
            {7'd73,7'd77}:		p = 14'd5621;
            {7'd73,7'd78}:		p = 14'd5694;
            {7'd73,7'd79}:		p = 14'd5767;
            {7'd73,7'd80}:		p = 14'd5840;
            {7'd73,7'd81}:		p = 14'd5913;
            {7'd73,7'd82}:		p = 14'd5986;
            {7'd73,7'd83}:		p = 14'd6059;
            {7'd73,7'd84}:		p = 14'd6132;
            {7'd73,7'd85}:		p = 14'd6205;
            {7'd73,7'd86}:		p = 14'd6278;
            {7'd73,7'd87}:		p = 14'd6351;
            {7'd73,7'd88}:		p = 14'd6424;
            {7'd73,7'd89}:		p = 14'd6497;
            {7'd73,7'd90}:		p = 14'd6570;
            {7'd73,7'd91}:		p = 14'd6643;
            {7'd73,7'd92}:		p = 14'd6716;
            {7'd73,7'd93}:		p = 14'd6789;
            {7'd73,7'd94}:		p = 14'd6862;
            {7'd73,7'd95}:		p = 14'd6935;
            {7'd73,7'd96}:		p = 14'd7008;
            {7'd73,7'd97}:		p = 14'd7081;
            {7'd73,7'd98}:		p = 14'd7154;
            {7'd73,7'd99}:		p = 14'd7227;
            {7'd73,7'd100}:		p = 14'd7300;
            {7'd73,7'd101}:		p = 14'd7373;
            {7'd73,7'd102}:		p = 14'd7446;
            {7'd73,7'd103}:		p = 14'd7519;
            {7'd73,7'd104}:		p = 14'd7592;
            {7'd73,7'd105}:		p = 14'd7665;
            {7'd73,7'd106}:		p = 14'd7738;
            {7'd73,7'd107}:		p = 14'd7811;
            {7'd73,7'd108}:		p = 14'd7884;
            {7'd73,7'd109}:		p = 14'd7957;
            {7'd73,7'd110}:		p = 14'd8030;
            {7'd73,7'd111}:		p = 14'd8103;
            {7'd73,7'd112}:		p = 14'd8176;
            {7'd73,7'd113}:		p = 14'd8249;
            {7'd73,7'd114}:		p = 14'd8322;
            {7'd73,7'd115}:		p = 14'd8395;
            {7'd73,7'd116}:		p = 14'd8468;
            {7'd73,7'd117}:		p = 14'd8541;
            {7'd73,7'd118}:		p = 14'd8614;
            {7'd73,7'd119}:		p = 14'd8687;
            {7'd73,7'd120}:		p = 14'd8760;
            {7'd73,7'd121}:		p = 14'd8833;
            {7'd73,7'd122}:		p = 14'd8906;
            {7'd73,7'd123}:		p = 14'd8979;
            {7'd73,7'd124}:		p = 14'd9052;
            {7'd73,7'd125}:		p = 14'd9125;
            {7'd73,7'd126}:		p = 14'd9198;
            {7'd73,7'd127}:		p = 14'd9271;
            {7'd74,7'd0}:		p = 14'd0;
            {7'd74,7'd1}:		p = 14'd74;
            {7'd74,7'd2}:		p = 14'd148;
            {7'd74,7'd3}:		p = 14'd222;
            {7'd74,7'd4}:		p = 14'd296;
            {7'd74,7'd5}:		p = 14'd370;
            {7'd74,7'd6}:		p = 14'd444;
            {7'd74,7'd7}:		p = 14'd518;
            {7'd74,7'd8}:		p = 14'd592;
            {7'd74,7'd9}:		p = 14'd666;
            {7'd74,7'd10}:		p = 14'd740;
            {7'd74,7'd11}:		p = 14'd814;
            {7'd74,7'd12}:		p = 14'd888;
            {7'd74,7'd13}:		p = 14'd962;
            {7'd74,7'd14}:		p = 14'd1036;
            {7'd74,7'd15}:		p = 14'd1110;
            {7'd74,7'd16}:		p = 14'd1184;
            {7'd74,7'd17}:		p = 14'd1258;
            {7'd74,7'd18}:		p = 14'd1332;
            {7'd74,7'd19}:		p = 14'd1406;
            {7'd74,7'd20}:		p = 14'd1480;
            {7'd74,7'd21}:		p = 14'd1554;
            {7'd74,7'd22}:		p = 14'd1628;
            {7'd74,7'd23}:		p = 14'd1702;
            {7'd74,7'd24}:		p = 14'd1776;
            {7'd74,7'd25}:		p = 14'd1850;
            {7'd74,7'd26}:		p = 14'd1924;
            {7'd74,7'd27}:		p = 14'd1998;
            {7'd74,7'd28}:		p = 14'd2072;
            {7'd74,7'd29}:		p = 14'd2146;
            {7'd74,7'd30}:		p = 14'd2220;
            {7'd74,7'd31}:		p = 14'd2294;
            {7'd74,7'd32}:		p = 14'd2368;
            {7'd74,7'd33}:		p = 14'd2442;
            {7'd74,7'd34}:		p = 14'd2516;
            {7'd74,7'd35}:		p = 14'd2590;
            {7'd74,7'd36}:		p = 14'd2664;
            {7'd74,7'd37}:		p = 14'd2738;
            {7'd74,7'd38}:		p = 14'd2812;
            {7'd74,7'd39}:		p = 14'd2886;
            {7'd74,7'd40}:		p = 14'd2960;
            {7'd74,7'd41}:		p = 14'd3034;
            {7'd74,7'd42}:		p = 14'd3108;
            {7'd74,7'd43}:		p = 14'd3182;
            {7'd74,7'd44}:		p = 14'd3256;
            {7'd74,7'd45}:		p = 14'd3330;
            {7'd74,7'd46}:		p = 14'd3404;
            {7'd74,7'd47}:		p = 14'd3478;
            {7'd74,7'd48}:		p = 14'd3552;
            {7'd74,7'd49}:		p = 14'd3626;
            {7'd74,7'd50}:		p = 14'd3700;
            {7'd74,7'd51}:		p = 14'd3774;
            {7'd74,7'd52}:		p = 14'd3848;
            {7'd74,7'd53}:		p = 14'd3922;
            {7'd74,7'd54}:		p = 14'd3996;
            {7'd74,7'd55}:		p = 14'd4070;
            {7'd74,7'd56}:		p = 14'd4144;
            {7'd74,7'd57}:		p = 14'd4218;
            {7'd74,7'd58}:		p = 14'd4292;
            {7'd74,7'd59}:		p = 14'd4366;
            {7'd74,7'd60}:		p = 14'd4440;
            {7'd74,7'd61}:		p = 14'd4514;
            {7'd74,7'd62}:		p = 14'd4588;
            {7'd74,7'd63}:		p = 14'd4662;
            {7'd74,7'd64}:		p = 14'd4736;
            {7'd74,7'd65}:		p = 14'd4810;
            {7'd74,7'd66}:		p = 14'd4884;
            {7'd74,7'd67}:		p = 14'd4958;
            {7'd74,7'd68}:		p = 14'd5032;
            {7'd74,7'd69}:		p = 14'd5106;
            {7'd74,7'd70}:		p = 14'd5180;
            {7'd74,7'd71}:		p = 14'd5254;
            {7'd74,7'd72}:		p = 14'd5328;
            {7'd74,7'd73}:		p = 14'd5402;
            {7'd74,7'd74}:		p = 14'd5476;
            {7'd74,7'd75}:		p = 14'd5550;
            {7'd74,7'd76}:		p = 14'd5624;
            {7'd74,7'd77}:		p = 14'd5698;
            {7'd74,7'd78}:		p = 14'd5772;
            {7'd74,7'd79}:		p = 14'd5846;
            {7'd74,7'd80}:		p = 14'd5920;
            {7'd74,7'd81}:		p = 14'd5994;
            {7'd74,7'd82}:		p = 14'd6068;
            {7'd74,7'd83}:		p = 14'd6142;
            {7'd74,7'd84}:		p = 14'd6216;
            {7'd74,7'd85}:		p = 14'd6290;
            {7'd74,7'd86}:		p = 14'd6364;
            {7'd74,7'd87}:		p = 14'd6438;
            {7'd74,7'd88}:		p = 14'd6512;
            {7'd74,7'd89}:		p = 14'd6586;
            {7'd74,7'd90}:		p = 14'd6660;
            {7'd74,7'd91}:		p = 14'd6734;
            {7'd74,7'd92}:		p = 14'd6808;
            {7'd74,7'd93}:		p = 14'd6882;
            {7'd74,7'd94}:		p = 14'd6956;
            {7'd74,7'd95}:		p = 14'd7030;
            {7'd74,7'd96}:		p = 14'd7104;
            {7'd74,7'd97}:		p = 14'd7178;
            {7'd74,7'd98}:		p = 14'd7252;
            {7'd74,7'd99}:		p = 14'd7326;
            {7'd74,7'd100}:		p = 14'd7400;
            {7'd74,7'd101}:		p = 14'd7474;
            {7'd74,7'd102}:		p = 14'd7548;
            {7'd74,7'd103}:		p = 14'd7622;
            {7'd74,7'd104}:		p = 14'd7696;
            {7'd74,7'd105}:		p = 14'd7770;
            {7'd74,7'd106}:		p = 14'd7844;
            {7'd74,7'd107}:		p = 14'd7918;
            {7'd74,7'd108}:		p = 14'd7992;
            {7'd74,7'd109}:		p = 14'd8066;
            {7'd74,7'd110}:		p = 14'd8140;
            {7'd74,7'd111}:		p = 14'd8214;
            {7'd74,7'd112}:		p = 14'd8288;
            {7'd74,7'd113}:		p = 14'd8362;
            {7'd74,7'd114}:		p = 14'd8436;
            {7'd74,7'd115}:		p = 14'd8510;
            {7'd74,7'd116}:		p = 14'd8584;
            {7'd74,7'd117}:		p = 14'd8658;
            {7'd74,7'd118}:		p = 14'd8732;
            {7'd74,7'd119}:		p = 14'd8806;
            {7'd74,7'd120}:		p = 14'd8880;
            {7'd74,7'd121}:		p = 14'd8954;
            {7'd74,7'd122}:		p = 14'd9028;
            {7'd74,7'd123}:		p = 14'd9102;
            {7'd74,7'd124}:		p = 14'd9176;
            {7'd74,7'd125}:		p = 14'd9250;
            {7'd74,7'd126}:		p = 14'd9324;
            {7'd74,7'd127}:		p = 14'd9398;
            {7'd75,7'd0}:		p = 14'd0;
            {7'd75,7'd1}:		p = 14'd75;
            {7'd75,7'd2}:		p = 14'd150;
            {7'd75,7'd3}:		p = 14'd225;
            {7'd75,7'd4}:		p = 14'd300;
            {7'd75,7'd5}:		p = 14'd375;
            {7'd75,7'd6}:		p = 14'd450;
            {7'd75,7'd7}:		p = 14'd525;
            {7'd75,7'd8}:		p = 14'd600;
            {7'd75,7'd9}:		p = 14'd675;
            {7'd75,7'd10}:		p = 14'd750;
            {7'd75,7'd11}:		p = 14'd825;
            {7'd75,7'd12}:		p = 14'd900;
            {7'd75,7'd13}:		p = 14'd975;
            {7'd75,7'd14}:		p = 14'd1050;
            {7'd75,7'd15}:		p = 14'd1125;
            {7'd75,7'd16}:		p = 14'd1200;
            {7'd75,7'd17}:		p = 14'd1275;
            {7'd75,7'd18}:		p = 14'd1350;
            {7'd75,7'd19}:		p = 14'd1425;
            {7'd75,7'd20}:		p = 14'd1500;
            {7'd75,7'd21}:		p = 14'd1575;
            {7'd75,7'd22}:		p = 14'd1650;
            {7'd75,7'd23}:		p = 14'd1725;
            {7'd75,7'd24}:		p = 14'd1800;
            {7'd75,7'd25}:		p = 14'd1875;
            {7'd75,7'd26}:		p = 14'd1950;
            {7'd75,7'd27}:		p = 14'd2025;
            {7'd75,7'd28}:		p = 14'd2100;
            {7'd75,7'd29}:		p = 14'd2175;
            {7'd75,7'd30}:		p = 14'd2250;
            {7'd75,7'd31}:		p = 14'd2325;
            {7'd75,7'd32}:		p = 14'd2400;
            {7'd75,7'd33}:		p = 14'd2475;
            {7'd75,7'd34}:		p = 14'd2550;
            {7'd75,7'd35}:		p = 14'd2625;
            {7'd75,7'd36}:		p = 14'd2700;
            {7'd75,7'd37}:		p = 14'd2775;
            {7'd75,7'd38}:		p = 14'd2850;
            {7'd75,7'd39}:		p = 14'd2925;
            {7'd75,7'd40}:		p = 14'd3000;
            {7'd75,7'd41}:		p = 14'd3075;
            {7'd75,7'd42}:		p = 14'd3150;
            {7'd75,7'd43}:		p = 14'd3225;
            {7'd75,7'd44}:		p = 14'd3300;
            {7'd75,7'd45}:		p = 14'd3375;
            {7'd75,7'd46}:		p = 14'd3450;
            {7'd75,7'd47}:		p = 14'd3525;
            {7'd75,7'd48}:		p = 14'd3600;
            {7'd75,7'd49}:		p = 14'd3675;
            {7'd75,7'd50}:		p = 14'd3750;
            {7'd75,7'd51}:		p = 14'd3825;
            {7'd75,7'd52}:		p = 14'd3900;
            {7'd75,7'd53}:		p = 14'd3975;
            {7'd75,7'd54}:		p = 14'd4050;
            {7'd75,7'd55}:		p = 14'd4125;
            {7'd75,7'd56}:		p = 14'd4200;
            {7'd75,7'd57}:		p = 14'd4275;
            {7'd75,7'd58}:		p = 14'd4350;
            {7'd75,7'd59}:		p = 14'd4425;
            {7'd75,7'd60}:		p = 14'd4500;
            {7'd75,7'd61}:		p = 14'd4575;
            {7'd75,7'd62}:		p = 14'd4650;
            {7'd75,7'd63}:		p = 14'd4725;
            {7'd75,7'd64}:		p = 14'd4800;
            {7'd75,7'd65}:		p = 14'd4875;
            {7'd75,7'd66}:		p = 14'd4950;
            {7'd75,7'd67}:		p = 14'd5025;
            {7'd75,7'd68}:		p = 14'd5100;
            {7'd75,7'd69}:		p = 14'd5175;
            {7'd75,7'd70}:		p = 14'd5250;
            {7'd75,7'd71}:		p = 14'd5325;
            {7'd75,7'd72}:		p = 14'd5400;
            {7'd75,7'd73}:		p = 14'd5475;
            {7'd75,7'd74}:		p = 14'd5550;
            {7'd75,7'd75}:		p = 14'd5625;
            {7'd75,7'd76}:		p = 14'd5700;
            {7'd75,7'd77}:		p = 14'd5775;
            {7'd75,7'd78}:		p = 14'd5850;
            {7'd75,7'd79}:		p = 14'd5925;
            {7'd75,7'd80}:		p = 14'd6000;
            {7'd75,7'd81}:		p = 14'd6075;
            {7'd75,7'd82}:		p = 14'd6150;
            {7'd75,7'd83}:		p = 14'd6225;
            {7'd75,7'd84}:		p = 14'd6300;
            {7'd75,7'd85}:		p = 14'd6375;
            {7'd75,7'd86}:		p = 14'd6450;
            {7'd75,7'd87}:		p = 14'd6525;
            {7'd75,7'd88}:		p = 14'd6600;
            {7'd75,7'd89}:		p = 14'd6675;
            {7'd75,7'd90}:		p = 14'd6750;
            {7'd75,7'd91}:		p = 14'd6825;
            {7'd75,7'd92}:		p = 14'd6900;
            {7'd75,7'd93}:		p = 14'd6975;
            {7'd75,7'd94}:		p = 14'd7050;
            {7'd75,7'd95}:		p = 14'd7125;
            {7'd75,7'd96}:		p = 14'd7200;
            {7'd75,7'd97}:		p = 14'd7275;
            {7'd75,7'd98}:		p = 14'd7350;
            {7'd75,7'd99}:		p = 14'd7425;
            {7'd75,7'd100}:		p = 14'd7500;
            {7'd75,7'd101}:		p = 14'd7575;
            {7'd75,7'd102}:		p = 14'd7650;
            {7'd75,7'd103}:		p = 14'd7725;
            {7'd75,7'd104}:		p = 14'd7800;
            {7'd75,7'd105}:		p = 14'd7875;
            {7'd75,7'd106}:		p = 14'd7950;
            {7'd75,7'd107}:		p = 14'd8025;
            {7'd75,7'd108}:		p = 14'd8100;
            {7'd75,7'd109}:		p = 14'd8175;
            {7'd75,7'd110}:		p = 14'd8250;
            {7'd75,7'd111}:		p = 14'd8325;
            {7'd75,7'd112}:		p = 14'd8400;
            {7'd75,7'd113}:		p = 14'd8475;
            {7'd75,7'd114}:		p = 14'd8550;
            {7'd75,7'd115}:		p = 14'd8625;
            {7'd75,7'd116}:		p = 14'd8700;
            {7'd75,7'd117}:		p = 14'd8775;
            {7'd75,7'd118}:		p = 14'd8850;
            {7'd75,7'd119}:		p = 14'd8925;
            {7'd75,7'd120}:		p = 14'd9000;
            {7'd75,7'd121}:		p = 14'd9075;
            {7'd75,7'd122}:		p = 14'd9150;
            {7'd75,7'd123}:		p = 14'd9225;
            {7'd75,7'd124}:		p = 14'd9300;
            {7'd75,7'd125}:		p = 14'd9375;
            {7'd75,7'd126}:		p = 14'd9450;
            {7'd75,7'd127}:		p = 14'd9525;
            {7'd76,7'd0}:		p = 14'd0;
            {7'd76,7'd1}:		p = 14'd76;
            {7'd76,7'd2}:		p = 14'd152;
            {7'd76,7'd3}:		p = 14'd228;
            {7'd76,7'd4}:		p = 14'd304;
            {7'd76,7'd5}:		p = 14'd380;
            {7'd76,7'd6}:		p = 14'd456;
            {7'd76,7'd7}:		p = 14'd532;
            {7'd76,7'd8}:		p = 14'd608;
            {7'd76,7'd9}:		p = 14'd684;
            {7'd76,7'd10}:		p = 14'd760;
            {7'd76,7'd11}:		p = 14'd836;
            {7'd76,7'd12}:		p = 14'd912;
            {7'd76,7'd13}:		p = 14'd988;
            {7'd76,7'd14}:		p = 14'd1064;
            {7'd76,7'd15}:		p = 14'd1140;
            {7'd76,7'd16}:		p = 14'd1216;
            {7'd76,7'd17}:		p = 14'd1292;
            {7'd76,7'd18}:		p = 14'd1368;
            {7'd76,7'd19}:		p = 14'd1444;
            {7'd76,7'd20}:		p = 14'd1520;
            {7'd76,7'd21}:		p = 14'd1596;
            {7'd76,7'd22}:		p = 14'd1672;
            {7'd76,7'd23}:		p = 14'd1748;
            {7'd76,7'd24}:		p = 14'd1824;
            {7'd76,7'd25}:		p = 14'd1900;
            {7'd76,7'd26}:		p = 14'd1976;
            {7'd76,7'd27}:		p = 14'd2052;
            {7'd76,7'd28}:		p = 14'd2128;
            {7'd76,7'd29}:		p = 14'd2204;
            {7'd76,7'd30}:		p = 14'd2280;
            {7'd76,7'd31}:		p = 14'd2356;
            {7'd76,7'd32}:		p = 14'd2432;
            {7'd76,7'd33}:		p = 14'd2508;
            {7'd76,7'd34}:		p = 14'd2584;
            {7'd76,7'd35}:		p = 14'd2660;
            {7'd76,7'd36}:		p = 14'd2736;
            {7'd76,7'd37}:		p = 14'd2812;
            {7'd76,7'd38}:		p = 14'd2888;
            {7'd76,7'd39}:		p = 14'd2964;
            {7'd76,7'd40}:		p = 14'd3040;
            {7'd76,7'd41}:		p = 14'd3116;
            {7'd76,7'd42}:		p = 14'd3192;
            {7'd76,7'd43}:		p = 14'd3268;
            {7'd76,7'd44}:		p = 14'd3344;
            {7'd76,7'd45}:		p = 14'd3420;
            {7'd76,7'd46}:		p = 14'd3496;
            {7'd76,7'd47}:		p = 14'd3572;
            {7'd76,7'd48}:		p = 14'd3648;
            {7'd76,7'd49}:		p = 14'd3724;
            {7'd76,7'd50}:		p = 14'd3800;
            {7'd76,7'd51}:		p = 14'd3876;
            {7'd76,7'd52}:		p = 14'd3952;
            {7'd76,7'd53}:		p = 14'd4028;
            {7'd76,7'd54}:		p = 14'd4104;
            {7'd76,7'd55}:		p = 14'd4180;
            {7'd76,7'd56}:		p = 14'd4256;
            {7'd76,7'd57}:		p = 14'd4332;
            {7'd76,7'd58}:		p = 14'd4408;
            {7'd76,7'd59}:		p = 14'd4484;
            {7'd76,7'd60}:		p = 14'd4560;
            {7'd76,7'd61}:		p = 14'd4636;
            {7'd76,7'd62}:		p = 14'd4712;
            {7'd76,7'd63}:		p = 14'd4788;
            {7'd76,7'd64}:		p = 14'd4864;
            {7'd76,7'd65}:		p = 14'd4940;
            {7'd76,7'd66}:		p = 14'd5016;
            {7'd76,7'd67}:		p = 14'd5092;
            {7'd76,7'd68}:		p = 14'd5168;
            {7'd76,7'd69}:		p = 14'd5244;
            {7'd76,7'd70}:		p = 14'd5320;
            {7'd76,7'd71}:		p = 14'd5396;
            {7'd76,7'd72}:		p = 14'd5472;
            {7'd76,7'd73}:		p = 14'd5548;
            {7'd76,7'd74}:		p = 14'd5624;
            {7'd76,7'd75}:		p = 14'd5700;
            {7'd76,7'd76}:		p = 14'd5776;
            {7'd76,7'd77}:		p = 14'd5852;
            {7'd76,7'd78}:		p = 14'd5928;
            {7'd76,7'd79}:		p = 14'd6004;
            {7'd76,7'd80}:		p = 14'd6080;
            {7'd76,7'd81}:		p = 14'd6156;
            {7'd76,7'd82}:		p = 14'd6232;
            {7'd76,7'd83}:		p = 14'd6308;
            {7'd76,7'd84}:		p = 14'd6384;
            {7'd76,7'd85}:		p = 14'd6460;
            {7'd76,7'd86}:		p = 14'd6536;
            {7'd76,7'd87}:		p = 14'd6612;
            {7'd76,7'd88}:		p = 14'd6688;
            {7'd76,7'd89}:		p = 14'd6764;
            {7'd76,7'd90}:		p = 14'd6840;
            {7'd76,7'd91}:		p = 14'd6916;
            {7'd76,7'd92}:		p = 14'd6992;
            {7'd76,7'd93}:		p = 14'd7068;
            {7'd76,7'd94}:		p = 14'd7144;
            {7'd76,7'd95}:		p = 14'd7220;
            {7'd76,7'd96}:		p = 14'd7296;
            {7'd76,7'd97}:		p = 14'd7372;
            {7'd76,7'd98}:		p = 14'd7448;
            {7'd76,7'd99}:		p = 14'd7524;
            {7'd76,7'd100}:		p = 14'd7600;
            {7'd76,7'd101}:		p = 14'd7676;
            {7'd76,7'd102}:		p = 14'd7752;
            {7'd76,7'd103}:		p = 14'd7828;
            {7'd76,7'd104}:		p = 14'd7904;
            {7'd76,7'd105}:		p = 14'd7980;
            {7'd76,7'd106}:		p = 14'd8056;
            {7'd76,7'd107}:		p = 14'd8132;
            {7'd76,7'd108}:		p = 14'd8208;
            {7'd76,7'd109}:		p = 14'd8284;
            {7'd76,7'd110}:		p = 14'd8360;
            {7'd76,7'd111}:		p = 14'd8436;
            {7'd76,7'd112}:		p = 14'd8512;
            {7'd76,7'd113}:		p = 14'd8588;
            {7'd76,7'd114}:		p = 14'd8664;
            {7'd76,7'd115}:		p = 14'd8740;
            {7'd76,7'd116}:		p = 14'd8816;
            {7'd76,7'd117}:		p = 14'd8892;
            {7'd76,7'd118}:		p = 14'd8968;
            {7'd76,7'd119}:		p = 14'd9044;
            {7'd76,7'd120}:		p = 14'd9120;
            {7'd76,7'd121}:		p = 14'd9196;
            {7'd76,7'd122}:		p = 14'd9272;
            {7'd76,7'd123}:		p = 14'd9348;
            {7'd76,7'd124}:		p = 14'd9424;
            {7'd76,7'd125}:		p = 14'd9500;
            {7'd76,7'd126}:		p = 14'd9576;
            {7'd76,7'd127}:		p = 14'd9652;
            {7'd77,7'd0}:		p = 14'd0;
            {7'd77,7'd1}:		p = 14'd77;
            {7'd77,7'd2}:		p = 14'd154;
            {7'd77,7'd3}:		p = 14'd231;
            {7'd77,7'd4}:		p = 14'd308;
            {7'd77,7'd5}:		p = 14'd385;
            {7'd77,7'd6}:		p = 14'd462;
            {7'd77,7'd7}:		p = 14'd539;
            {7'd77,7'd8}:		p = 14'd616;
            {7'd77,7'd9}:		p = 14'd693;
            {7'd77,7'd10}:		p = 14'd770;
            {7'd77,7'd11}:		p = 14'd847;
            {7'd77,7'd12}:		p = 14'd924;
            {7'd77,7'd13}:		p = 14'd1001;
            {7'd77,7'd14}:		p = 14'd1078;
            {7'd77,7'd15}:		p = 14'd1155;
            {7'd77,7'd16}:		p = 14'd1232;
            {7'd77,7'd17}:		p = 14'd1309;
            {7'd77,7'd18}:		p = 14'd1386;
            {7'd77,7'd19}:		p = 14'd1463;
            {7'd77,7'd20}:		p = 14'd1540;
            {7'd77,7'd21}:		p = 14'd1617;
            {7'd77,7'd22}:		p = 14'd1694;
            {7'd77,7'd23}:		p = 14'd1771;
            {7'd77,7'd24}:		p = 14'd1848;
            {7'd77,7'd25}:		p = 14'd1925;
            {7'd77,7'd26}:		p = 14'd2002;
            {7'd77,7'd27}:		p = 14'd2079;
            {7'd77,7'd28}:		p = 14'd2156;
            {7'd77,7'd29}:		p = 14'd2233;
            {7'd77,7'd30}:		p = 14'd2310;
            {7'd77,7'd31}:		p = 14'd2387;
            {7'd77,7'd32}:		p = 14'd2464;
            {7'd77,7'd33}:		p = 14'd2541;
            {7'd77,7'd34}:		p = 14'd2618;
            {7'd77,7'd35}:		p = 14'd2695;
            {7'd77,7'd36}:		p = 14'd2772;
            {7'd77,7'd37}:		p = 14'd2849;
            {7'd77,7'd38}:		p = 14'd2926;
            {7'd77,7'd39}:		p = 14'd3003;
            {7'd77,7'd40}:		p = 14'd3080;
            {7'd77,7'd41}:		p = 14'd3157;
            {7'd77,7'd42}:		p = 14'd3234;
            {7'd77,7'd43}:		p = 14'd3311;
            {7'd77,7'd44}:		p = 14'd3388;
            {7'd77,7'd45}:		p = 14'd3465;
            {7'd77,7'd46}:		p = 14'd3542;
            {7'd77,7'd47}:		p = 14'd3619;
            {7'd77,7'd48}:		p = 14'd3696;
            {7'd77,7'd49}:		p = 14'd3773;
            {7'd77,7'd50}:		p = 14'd3850;
            {7'd77,7'd51}:		p = 14'd3927;
            {7'd77,7'd52}:		p = 14'd4004;
            {7'd77,7'd53}:		p = 14'd4081;
            {7'd77,7'd54}:		p = 14'd4158;
            {7'd77,7'd55}:		p = 14'd4235;
            {7'd77,7'd56}:		p = 14'd4312;
            {7'd77,7'd57}:		p = 14'd4389;
            {7'd77,7'd58}:		p = 14'd4466;
            {7'd77,7'd59}:		p = 14'd4543;
            {7'd77,7'd60}:		p = 14'd4620;
            {7'd77,7'd61}:		p = 14'd4697;
            {7'd77,7'd62}:		p = 14'd4774;
            {7'd77,7'd63}:		p = 14'd4851;
            {7'd77,7'd64}:		p = 14'd4928;
            {7'd77,7'd65}:		p = 14'd5005;
            {7'd77,7'd66}:		p = 14'd5082;
            {7'd77,7'd67}:		p = 14'd5159;
            {7'd77,7'd68}:		p = 14'd5236;
            {7'd77,7'd69}:		p = 14'd5313;
            {7'd77,7'd70}:		p = 14'd5390;
            {7'd77,7'd71}:		p = 14'd5467;
            {7'd77,7'd72}:		p = 14'd5544;
            {7'd77,7'd73}:		p = 14'd5621;
            {7'd77,7'd74}:		p = 14'd5698;
            {7'd77,7'd75}:		p = 14'd5775;
            {7'd77,7'd76}:		p = 14'd5852;
            {7'd77,7'd77}:		p = 14'd5929;
            {7'd77,7'd78}:		p = 14'd6006;
            {7'd77,7'd79}:		p = 14'd6083;
            {7'd77,7'd80}:		p = 14'd6160;
            {7'd77,7'd81}:		p = 14'd6237;
            {7'd77,7'd82}:		p = 14'd6314;
            {7'd77,7'd83}:		p = 14'd6391;
            {7'd77,7'd84}:		p = 14'd6468;
            {7'd77,7'd85}:		p = 14'd6545;
            {7'd77,7'd86}:		p = 14'd6622;
            {7'd77,7'd87}:		p = 14'd6699;
            {7'd77,7'd88}:		p = 14'd6776;
            {7'd77,7'd89}:		p = 14'd6853;
            {7'd77,7'd90}:		p = 14'd6930;
            {7'd77,7'd91}:		p = 14'd7007;
            {7'd77,7'd92}:		p = 14'd7084;
            {7'd77,7'd93}:		p = 14'd7161;
            {7'd77,7'd94}:		p = 14'd7238;
            {7'd77,7'd95}:		p = 14'd7315;
            {7'd77,7'd96}:		p = 14'd7392;
            {7'd77,7'd97}:		p = 14'd7469;
            {7'd77,7'd98}:		p = 14'd7546;
            {7'd77,7'd99}:		p = 14'd7623;
            {7'd77,7'd100}:		p = 14'd7700;
            {7'd77,7'd101}:		p = 14'd7777;
            {7'd77,7'd102}:		p = 14'd7854;
            {7'd77,7'd103}:		p = 14'd7931;
            {7'd77,7'd104}:		p = 14'd8008;
            {7'd77,7'd105}:		p = 14'd8085;
            {7'd77,7'd106}:		p = 14'd8162;
            {7'd77,7'd107}:		p = 14'd8239;
            {7'd77,7'd108}:		p = 14'd8316;
            {7'd77,7'd109}:		p = 14'd8393;
            {7'd77,7'd110}:		p = 14'd8470;
            {7'd77,7'd111}:		p = 14'd8547;
            {7'd77,7'd112}:		p = 14'd8624;
            {7'd77,7'd113}:		p = 14'd8701;
            {7'd77,7'd114}:		p = 14'd8778;
            {7'd77,7'd115}:		p = 14'd8855;
            {7'd77,7'd116}:		p = 14'd8932;
            {7'd77,7'd117}:		p = 14'd9009;
            {7'd77,7'd118}:		p = 14'd9086;
            {7'd77,7'd119}:		p = 14'd9163;
            {7'd77,7'd120}:		p = 14'd9240;
            {7'd77,7'd121}:		p = 14'd9317;
            {7'd77,7'd122}:		p = 14'd9394;
            {7'd77,7'd123}:		p = 14'd9471;
            {7'd77,7'd124}:		p = 14'd9548;
            {7'd77,7'd125}:		p = 14'd9625;
            {7'd77,7'd126}:		p = 14'd9702;
            {7'd77,7'd127}:		p = 14'd9779;
            {7'd78,7'd0}:		p = 14'd0;
            {7'd78,7'd1}:		p = 14'd78;
            {7'd78,7'd2}:		p = 14'd156;
            {7'd78,7'd3}:		p = 14'd234;
            {7'd78,7'd4}:		p = 14'd312;
            {7'd78,7'd5}:		p = 14'd390;
            {7'd78,7'd6}:		p = 14'd468;
            {7'd78,7'd7}:		p = 14'd546;
            {7'd78,7'd8}:		p = 14'd624;
            {7'd78,7'd9}:		p = 14'd702;
            {7'd78,7'd10}:		p = 14'd780;
            {7'd78,7'd11}:		p = 14'd858;
            {7'd78,7'd12}:		p = 14'd936;
            {7'd78,7'd13}:		p = 14'd1014;
            {7'd78,7'd14}:		p = 14'd1092;
            {7'd78,7'd15}:		p = 14'd1170;
            {7'd78,7'd16}:		p = 14'd1248;
            {7'd78,7'd17}:		p = 14'd1326;
            {7'd78,7'd18}:		p = 14'd1404;
            {7'd78,7'd19}:		p = 14'd1482;
            {7'd78,7'd20}:		p = 14'd1560;
            {7'd78,7'd21}:		p = 14'd1638;
            {7'd78,7'd22}:		p = 14'd1716;
            {7'd78,7'd23}:		p = 14'd1794;
            {7'd78,7'd24}:		p = 14'd1872;
            {7'd78,7'd25}:		p = 14'd1950;
            {7'd78,7'd26}:		p = 14'd2028;
            {7'd78,7'd27}:		p = 14'd2106;
            {7'd78,7'd28}:		p = 14'd2184;
            {7'd78,7'd29}:		p = 14'd2262;
            {7'd78,7'd30}:		p = 14'd2340;
            {7'd78,7'd31}:		p = 14'd2418;
            {7'd78,7'd32}:		p = 14'd2496;
            {7'd78,7'd33}:		p = 14'd2574;
            {7'd78,7'd34}:		p = 14'd2652;
            {7'd78,7'd35}:		p = 14'd2730;
            {7'd78,7'd36}:		p = 14'd2808;
            {7'd78,7'd37}:		p = 14'd2886;
            {7'd78,7'd38}:		p = 14'd2964;
            {7'd78,7'd39}:		p = 14'd3042;
            {7'd78,7'd40}:		p = 14'd3120;
            {7'd78,7'd41}:		p = 14'd3198;
            {7'd78,7'd42}:		p = 14'd3276;
            {7'd78,7'd43}:		p = 14'd3354;
            {7'd78,7'd44}:		p = 14'd3432;
            {7'd78,7'd45}:		p = 14'd3510;
            {7'd78,7'd46}:		p = 14'd3588;
            {7'd78,7'd47}:		p = 14'd3666;
            {7'd78,7'd48}:		p = 14'd3744;
            {7'd78,7'd49}:		p = 14'd3822;
            {7'd78,7'd50}:		p = 14'd3900;
            {7'd78,7'd51}:		p = 14'd3978;
            {7'd78,7'd52}:		p = 14'd4056;
            {7'd78,7'd53}:		p = 14'd4134;
            {7'd78,7'd54}:		p = 14'd4212;
            {7'd78,7'd55}:		p = 14'd4290;
            {7'd78,7'd56}:		p = 14'd4368;
            {7'd78,7'd57}:		p = 14'd4446;
            {7'd78,7'd58}:		p = 14'd4524;
            {7'd78,7'd59}:		p = 14'd4602;
            {7'd78,7'd60}:		p = 14'd4680;
            {7'd78,7'd61}:		p = 14'd4758;
            {7'd78,7'd62}:		p = 14'd4836;
            {7'd78,7'd63}:		p = 14'd4914;
            {7'd78,7'd64}:		p = 14'd4992;
            {7'd78,7'd65}:		p = 14'd5070;
            {7'd78,7'd66}:		p = 14'd5148;
            {7'd78,7'd67}:		p = 14'd5226;
            {7'd78,7'd68}:		p = 14'd5304;
            {7'd78,7'd69}:		p = 14'd5382;
            {7'd78,7'd70}:		p = 14'd5460;
            {7'd78,7'd71}:		p = 14'd5538;
            {7'd78,7'd72}:		p = 14'd5616;
            {7'd78,7'd73}:		p = 14'd5694;
            {7'd78,7'd74}:		p = 14'd5772;
            {7'd78,7'd75}:		p = 14'd5850;
            {7'd78,7'd76}:		p = 14'd5928;
            {7'd78,7'd77}:		p = 14'd6006;
            {7'd78,7'd78}:		p = 14'd6084;
            {7'd78,7'd79}:		p = 14'd6162;
            {7'd78,7'd80}:		p = 14'd6240;
            {7'd78,7'd81}:		p = 14'd6318;
            {7'd78,7'd82}:		p = 14'd6396;
            {7'd78,7'd83}:		p = 14'd6474;
            {7'd78,7'd84}:		p = 14'd6552;
            {7'd78,7'd85}:		p = 14'd6630;
            {7'd78,7'd86}:		p = 14'd6708;
            {7'd78,7'd87}:		p = 14'd6786;
            {7'd78,7'd88}:		p = 14'd6864;
            {7'd78,7'd89}:		p = 14'd6942;
            {7'd78,7'd90}:		p = 14'd7020;
            {7'd78,7'd91}:		p = 14'd7098;
            {7'd78,7'd92}:		p = 14'd7176;
            {7'd78,7'd93}:		p = 14'd7254;
            {7'd78,7'd94}:		p = 14'd7332;
            {7'd78,7'd95}:		p = 14'd7410;
            {7'd78,7'd96}:		p = 14'd7488;
            {7'd78,7'd97}:		p = 14'd7566;
            {7'd78,7'd98}:		p = 14'd7644;
            {7'd78,7'd99}:		p = 14'd7722;
            {7'd78,7'd100}:		p = 14'd7800;
            {7'd78,7'd101}:		p = 14'd7878;
            {7'd78,7'd102}:		p = 14'd7956;
            {7'd78,7'd103}:		p = 14'd8034;
            {7'd78,7'd104}:		p = 14'd8112;
            {7'd78,7'd105}:		p = 14'd8190;
            {7'd78,7'd106}:		p = 14'd8268;
            {7'd78,7'd107}:		p = 14'd8346;
            {7'd78,7'd108}:		p = 14'd8424;
            {7'd78,7'd109}:		p = 14'd8502;
            {7'd78,7'd110}:		p = 14'd8580;
            {7'd78,7'd111}:		p = 14'd8658;
            {7'd78,7'd112}:		p = 14'd8736;
            {7'd78,7'd113}:		p = 14'd8814;
            {7'd78,7'd114}:		p = 14'd8892;
            {7'd78,7'd115}:		p = 14'd8970;
            {7'd78,7'd116}:		p = 14'd9048;
            {7'd78,7'd117}:		p = 14'd9126;
            {7'd78,7'd118}:		p = 14'd9204;
            {7'd78,7'd119}:		p = 14'd9282;
            {7'd78,7'd120}:		p = 14'd9360;
            {7'd78,7'd121}:		p = 14'd9438;
            {7'd78,7'd122}:		p = 14'd9516;
            {7'd78,7'd123}:		p = 14'd9594;
            {7'd78,7'd124}:		p = 14'd9672;
            {7'd78,7'd125}:		p = 14'd9750;
            {7'd78,7'd126}:		p = 14'd9828;
            {7'd78,7'd127}:		p = 14'd9906;
            {7'd79,7'd0}:		p = 14'd0;
            {7'd79,7'd1}:		p = 14'd79;
            {7'd79,7'd2}:		p = 14'd158;
            {7'd79,7'd3}:		p = 14'd237;
            {7'd79,7'd4}:		p = 14'd316;
            {7'd79,7'd5}:		p = 14'd395;
            {7'd79,7'd6}:		p = 14'd474;
            {7'd79,7'd7}:		p = 14'd553;
            {7'd79,7'd8}:		p = 14'd632;
            {7'd79,7'd9}:		p = 14'd711;
            {7'd79,7'd10}:		p = 14'd790;
            {7'd79,7'd11}:		p = 14'd869;
            {7'd79,7'd12}:		p = 14'd948;
            {7'd79,7'd13}:		p = 14'd1027;
            {7'd79,7'd14}:		p = 14'd1106;
            {7'd79,7'd15}:		p = 14'd1185;
            {7'd79,7'd16}:		p = 14'd1264;
            {7'd79,7'd17}:		p = 14'd1343;
            {7'd79,7'd18}:		p = 14'd1422;
            {7'd79,7'd19}:		p = 14'd1501;
            {7'd79,7'd20}:		p = 14'd1580;
            {7'd79,7'd21}:		p = 14'd1659;
            {7'd79,7'd22}:		p = 14'd1738;
            {7'd79,7'd23}:		p = 14'd1817;
            {7'd79,7'd24}:		p = 14'd1896;
            {7'd79,7'd25}:		p = 14'd1975;
            {7'd79,7'd26}:		p = 14'd2054;
            {7'd79,7'd27}:		p = 14'd2133;
            {7'd79,7'd28}:		p = 14'd2212;
            {7'd79,7'd29}:		p = 14'd2291;
            {7'd79,7'd30}:		p = 14'd2370;
            {7'd79,7'd31}:		p = 14'd2449;
            {7'd79,7'd32}:		p = 14'd2528;
            {7'd79,7'd33}:		p = 14'd2607;
            {7'd79,7'd34}:		p = 14'd2686;
            {7'd79,7'd35}:		p = 14'd2765;
            {7'd79,7'd36}:		p = 14'd2844;
            {7'd79,7'd37}:		p = 14'd2923;
            {7'd79,7'd38}:		p = 14'd3002;
            {7'd79,7'd39}:		p = 14'd3081;
            {7'd79,7'd40}:		p = 14'd3160;
            {7'd79,7'd41}:		p = 14'd3239;
            {7'd79,7'd42}:		p = 14'd3318;
            {7'd79,7'd43}:		p = 14'd3397;
            {7'd79,7'd44}:		p = 14'd3476;
            {7'd79,7'd45}:		p = 14'd3555;
            {7'd79,7'd46}:		p = 14'd3634;
            {7'd79,7'd47}:		p = 14'd3713;
            {7'd79,7'd48}:		p = 14'd3792;
            {7'd79,7'd49}:		p = 14'd3871;
            {7'd79,7'd50}:		p = 14'd3950;
            {7'd79,7'd51}:		p = 14'd4029;
            {7'd79,7'd52}:		p = 14'd4108;
            {7'd79,7'd53}:		p = 14'd4187;
            {7'd79,7'd54}:		p = 14'd4266;
            {7'd79,7'd55}:		p = 14'd4345;
            {7'd79,7'd56}:		p = 14'd4424;
            {7'd79,7'd57}:		p = 14'd4503;
            {7'd79,7'd58}:		p = 14'd4582;
            {7'd79,7'd59}:		p = 14'd4661;
            {7'd79,7'd60}:		p = 14'd4740;
            {7'd79,7'd61}:		p = 14'd4819;
            {7'd79,7'd62}:		p = 14'd4898;
            {7'd79,7'd63}:		p = 14'd4977;
            {7'd79,7'd64}:		p = 14'd5056;
            {7'd79,7'd65}:		p = 14'd5135;
            {7'd79,7'd66}:		p = 14'd5214;
            {7'd79,7'd67}:		p = 14'd5293;
            {7'd79,7'd68}:		p = 14'd5372;
            {7'd79,7'd69}:		p = 14'd5451;
            {7'd79,7'd70}:		p = 14'd5530;
            {7'd79,7'd71}:		p = 14'd5609;
            {7'd79,7'd72}:		p = 14'd5688;
            {7'd79,7'd73}:		p = 14'd5767;
            {7'd79,7'd74}:		p = 14'd5846;
            {7'd79,7'd75}:		p = 14'd5925;
            {7'd79,7'd76}:		p = 14'd6004;
            {7'd79,7'd77}:		p = 14'd6083;
            {7'd79,7'd78}:		p = 14'd6162;
            {7'd79,7'd79}:		p = 14'd6241;
            {7'd79,7'd80}:		p = 14'd6320;
            {7'd79,7'd81}:		p = 14'd6399;
            {7'd79,7'd82}:		p = 14'd6478;
            {7'd79,7'd83}:		p = 14'd6557;
            {7'd79,7'd84}:		p = 14'd6636;
            {7'd79,7'd85}:		p = 14'd6715;
            {7'd79,7'd86}:		p = 14'd6794;
            {7'd79,7'd87}:		p = 14'd6873;
            {7'd79,7'd88}:		p = 14'd6952;
            {7'd79,7'd89}:		p = 14'd7031;
            {7'd79,7'd90}:		p = 14'd7110;
            {7'd79,7'd91}:		p = 14'd7189;
            {7'd79,7'd92}:		p = 14'd7268;
            {7'd79,7'd93}:		p = 14'd7347;
            {7'd79,7'd94}:		p = 14'd7426;
            {7'd79,7'd95}:		p = 14'd7505;
            {7'd79,7'd96}:		p = 14'd7584;
            {7'd79,7'd97}:		p = 14'd7663;
            {7'd79,7'd98}:		p = 14'd7742;
            {7'd79,7'd99}:		p = 14'd7821;
            {7'd79,7'd100}:		p = 14'd7900;
            {7'd79,7'd101}:		p = 14'd7979;
            {7'd79,7'd102}:		p = 14'd8058;
            {7'd79,7'd103}:		p = 14'd8137;
            {7'd79,7'd104}:		p = 14'd8216;
            {7'd79,7'd105}:		p = 14'd8295;
            {7'd79,7'd106}:		p = 14'd8374;
            {7'd79,7'd107}:		p = 14'd8453;
            {7'd79,7'd108}:		p = 14'd8532;
            {7'd79,7'd109}:		p = 14'd8611;
            {7'd79,7'd110}:		p = 14'd8690;
            {7'd79,7'd111}:		p = 14'd8769;
            {7'd79,7'd112}:		p = 14'd8848;
            {7'd79,7'd113}:		p = 14'd8927;
            {7'd79,7'd114}:		p = 14'd9006;
            {7'd79,7'd115}:		p = 14'd9085;
            {7'd79,7'd116}:		p = 14'd9164;
            {7'd79,7'd117}:		p = 14'd9243;
            {7'd79,7'd118}:		p = 14'd9322;
            {7'd79,7'd119}:		p = 14'd9401;
            {7'd79,7'd120}:		p = 14'd9480;
            {7'd79,7'd121}:		p = 14'd9559;
            {7'd79,7'd122}:		p = 14'd9638;
            {7'd79,7'd123}:		p = 14'd9717;
            {7'd79,7'd124}:		p = 14'd9796;
            {7'd79,7'd125}:		p = 14'd9875;
            {7'd79,7'd126}:		p = 14'd9954;
            {7'd79,7'd127}:		p = 14'd10033;
            {7'd80,7'd0}:		p = 14'd0;
            {7'd80,7'd1}:		p = 14'd80;
            {7'd80,7'd2}:		p = 14'd160;
            {7'd80,7'd3}:		p = 14'd240;
            {7'd80,7'd4}:		p = 14'd320;
            {7'd80,7'd5}:		p = 14'd400;
            {7'd80,7'd6}:		p = 14'd480;
            {7'd80,7'd7}:		p = 14'd560;
            {7'd80,7'd8}:		p = 14'd640;
            {7'd80,7'd9}:		p = 14'd720;
            {7'd80,7'd10}:		p = 14'd800;
            {7'd80,7'd11}:		p = 14'd880;
            {7'd80,7'd12}:		p = 14'd960;
            {7'd80,7'd13}:		p = 14'd1040;
            {7'd80,7'd14}:		p = 14'd1120;
            {7'd80,7'd15}:		p = 14'd1200;
            {7'd80,7'd16}:		p = 14'd1280;
            {7'd80,7'd17}:		p = 14'd1360;
            {7'd80,7'd18}:		p = 14'd1440;
            {7'd80,7'd19}:		p = 14'd1520;
            {7'd80,7'd20}:		p = 14'd1600;
            {7'd80,7'd21}:		p = 14'd1680;
            {7'd80,7'd22}:		p = 14'd1760;
            {7'd80,7'd23}:		p = 14'd1840;
            {7'd80,7'd24}:		p = 14'd1920;
            {7'd80,7'd25}:		p = 14'd2000;
            {7'd80,7'd26}:		p = 14'd2080;
            {7'd80,7'd27}:		p = 14'd2160;
            {7'd80,7'd28}:		p = 14'd2240;
            {7'd80,7'd29}:		p = 14'd2320;
            {7'd80,7'd30}:		p = 14'd2400;
            {7'd80,7'd31}:		p = 14'd2480;
            {7'd80,7'd32}:		p = 14'd2560;
            {7'd80,7'd33}:		p = 14'd2640;
            {7'd80,7'd34}:		p = 14'd2720;
            {7'd80,7'd35}:		p = 14'd2800;
            {7'd80,7'd36}:		p = 14'd2880;
            {7'd80,7'd37}:		p = 14'd2960;
            {7'd80,7'd38}:		p = 14'd3040;
            {7'd80,7'd39}:		p = 14'd3120;
            {7'd80,7'd40}:		p = 14'd3200;
            {7'd80,7'd41}:		p = 14'd3280;
            {7'd80,7'd42}:		p = 14'd3360;
            {7'd80,7'd43}:		p = 14'd3440;
            {7'd80,7'd44}:		p = 14'd3520;
            {7'd80,7'd45}:		p = 14'd3600;
            {7'd80,7'd46}:		p = 14'd3680;
            {7'd80,7'd47}:		p = 14'd3760;
            {7'd80,7'd48}:		p = 14'd3840;
            {7'd80,7'd49}:		p = 14'd3920;
            {7'd80,7'd50}:		p = 14'd4000;
            {7'd80,7'd51}:		p = 14'd4080;
            {7'd80,7'd52}:		p = 14'd4160;
            {7'd80,7'd53}:		p = 14'd4240;
            {7'd80,7'd54}:		p = 14'd4320;
            {7'd80,7'd55}:		p = 14'd4400;
            {7'd80,7'd56}:		p = 14'd4480;
            {7'd80,7'd57}:		p = 14'd4560;
            {7'd80,7'd58}:		p = 14'd4640;
            {7'd80,7'd59}:		p = 14'd4720;
            {7'd80,7'd60}:		p = 14'd4800;
            {7'd80,7'd61}:		p = 14'd4880;
            {7'd80,7'd62}:		p = 14'd4960;
            {7'd80,7'd63}:		p = 14'd5040;
            {7'd80,7'd64}:		p = 14'd5120;
            {7'd80,7'd65}:		p = 14'd5200;
            {7'd80,7'd66}:		p = 14'd5280;
            {7'd80,7'd67}:		p = 14'd5360;
            {7'd80,7'd68}:		p = 14'd5440;
            {7'd80,7'd69}:		p = 14'd5520;
            {7'd80,7'd70}:		p = 14'd5600;
            {7'd80,7'd71}:		p = 14'd5680;
            {7'd80,7'd72}:		p = 14'd5760;
            {7'd80,7'd73}:		p = 14'd5840;
            {7'd80,7'd74}:		p = 14'd5920;
            {7'd80,7'd75}:		p = 14'd6000;
            {7'd80,7'd76}:		p = 14'd6080;
            {7'd80,7'd77}:		p = 14'd6160;
            {7'd80,7'd78}:		p = 14'd6240;
            {7'd80,7'd79}:		p = 14'd6320;
            {7'd80,7'd80}:		p = 14'd6400;
            {7'd80,7'd81}:		p = 14'd6480;
            {7'd80,7'd82}:		p = 14'd6560;
            {7'd80,7'd83}:		p = 14'd6640;
            {7'd80,7'd84}:		p = 14'd6720;
            {7'd80,7'd85}:		p = 14'd6800;
            {7'd80,7'd86}:		p = 14'd6880;
            {7'd80,7'd87}:		p = 14'd6960;
            {7'd80,7'd88}:		p = 14'd7040;
            {7'd80,7'd89}:		p = 14'd7120;
            {7'd80,7'd90}:		p = 14'd7200;
            {7'd80,7'd91}:		p = 14'd7280;
            {7'd80,7'd92}:		p = 14'd7360;
            {7'd80,7'd93}:		p = 14'd7440;
            {7'd80,7'd94}:		p = 14'd7520;
            {7'd80,7'd95}:		p = 14'd7600;
            {7'd80,7'd96}:		p = 14'd7680;
            {7'd80,7'd97}:		p = 14'd7760;
            {7'd80,7'd98}:		p = 14'd7840;
            {7'd80,7'd99}:		p = 14'd7920;
            {7'd80,7'd100}:		p = 14'd8000;
            {7'd80,7'd101}:		p = 14'd8080;
            {7'd80,7'd102}:		p = 14'd8160;
            {7'd80,7'd103}:		p = 14'd8240;
            {7'd80,7'd104}:		p = 14'd8320;
            {7'd80,7'd105}:		p = 14'd8400;
            {7'd80,7'd106}:		p = 14'd8480;
            {7'd80,7'd107}:		p = 14'd8560;
            {7'd80,7'd108}:		p = 14'd8640;
            {7'd80,7'd109}:		p = 14'd8720;
            {7'd80,7'd110}:		p = 14'd8800;
            {7'd80,7'd111}:		p = 14'd8880;
            {7'd80,7'd112}:		p = 14'd8960;
            {7'd80,7'd113}:		p = 14'd9040;
            {7'd80,7'd114}:		p = 14'd9120;
            {7'd80,7'd115}:		p = 14'd9200;
            {7'd80,7'd116}:		p = 14'd9280;
            {7'd80,7'd117}:		p = 14'd9360;
            {7'd80,7'd118}:		p = 14'd9440;
            {7'd80,7'd119}:		p = 14'd9520;
            {7'd80,7'd120}:		p = 14'd9600;
            {7'd80,7'd121}:		p = 14'd9680;
            {7'd80,7'd122}:		p = 14'd9760;
            {7'd80,7'd123}:		p = 14'd9840;
            {7'd80,7'd124}:		p = 14'd9920;
            {7'd80,7'd125}:		p = 14'd10000;
            {7'd80,7'd126}:		p = 14'd10080;
            {7'd80,7'd127}:		p = 14'd10160;
            {7'd81,7'd0}:		p = 14'd0;
            {7'd81,7'd1}:		p = 14'd81;
            {7'd81,7'd2}:		p = 14'd162;
            {7'd81,7'd3}:		p = 14'd243;
            {7'd81,7'd4}:		p = 14'd324;
            {7'd81,7'd5}:		p = 14'd405;
            {7'd81,7'd6}:		p = 14'd486;
            {7'd81,7'd7}:		p = 14'd567;
            {7'd81,7'd8}:		p = 14'd648;
            {7'd81,7'd9}:		p = 14'd729;
            {7'd81,7'd10}:		p = 14'd810;
            {7'd81,7'd11}:		p = 14'd891;
            {7'd81,7'd12}:		p = 14'd972;
            {7'd81,7'd13}:		p = 14'd1053;
            {7'd81,7'd14}:		p = 14'd1134;
            {7'd81,7'd15}:		p = 14'd1215;
            {7'd81,7'd16}:		p = 14'd1296;
            {7'd81,7'd17}:		p = 14'd1377;
            {7'd81,7'd18}:		p = 14'd1458;
            {7'd81,7'd19}:		p = 14'd1539;
            {7'd81,7'd20}:		p = 14'd1620;
            {7'd81,7'd21}:		p = 14'd1701;
            {7'd81,7'd22}:		p = 14'd1782;
            {7'd81,7'd23}:		p = 14'd1863;
            {7'd81,7'd24}:		p = 14'd1944;
            {7'd81,7'd25}:		p = 14'd2025;
            {7'd81,7'd26}:		p = 14'd2106;
            {7'd81,7'd27}:		p = 14'd2187;
            {7'd81,7'd28}:		p = 14'd2268;
            {7'd81,7'd29}:		p = 14'd2349;
            {7'd81,7'd30}:		p = 14'd2430;
            {7'd81,7'd31}:		p = 14'd2511;
            {7'd81,7'd32}:		p = 14'd2592;
            {7'd81,7'd33}:		p = 14'd2673;
            {7'd81,7'd34}:		p = 14'd2754;
            {7'd81,7'd35}:		p = 14'd2835;
            {7'd81,7'd36}:		p = 14'd2916;
            {7'd81,7'd37}:		p = 14'd2997;
            {7'd81,7'd38}:		p = 14'd3078;
            {7'd81,7'd39}:		p = 14'd3159;
            {7'd81,7'd40}:		p = 14'd3240;
            {7'd81,7'd41}:		p = 14'd3321;
            {7'd81,7'd42}:		p = 14'd3402;
            {7'd81,7'd43}:		p = 14'd3483;
            {7'd81,7'd44}:		p = 14'd3564;
            {7'd81,7'd45}:		p = 14'd3645;
            {7'd81,7'd46}:		p = 14'd3726;
            {7'd81,7'd47}:		p = 14'd3807;
            {7'd81,7'd48}:		p = 14'd3888;
            {7'd81,7'd49}:		p = 14'd3969;
            {7'd81,7'd50}:		p = 14'd4050;
            {7'd81,7'd51}:		p = 14'd4131;
            {7'd81,7'd52}:		p = 14'd4212;
            {7'd81,7'd53}:		p = 14'd4293;
            {7'd81,7'd54}:		p = 14'd4374;
            {7'd81,7'd55}:		p = 14'd4455;
            {7'd81,7'd56}:		p = 14'd4536;
            {7'd81,7'd57}:		p = 14'd4617;
            {7'd81,7'd58}:		p = 14'd4698;
            {7'd81,7'd59}:		p = 14'd4779;
            {7'd81,7'd60}:		p = 14'd4860;
            {7'd81,7'd61}:		p = 14'd4941;
            {7'd81,7'd62}:		p = 14'd5022;
            {7'd81,7'd63}:		p = 14'd5103;
            {7'd81,7'd64}:		p = 14'd5184;
            {7'd81,7'd65}:		p = 14'd5265;
            {7'd81,7'd66}:		p = 14'd5346;
            {7'd81,7'd67}:		p = 14'd5427;
            {7'd81,7'd68}:		p = 14'd5508;
            {7'd81,7'd69}:		p = 14'd5589;
            {7'd81,7'd70}:		p = 14'd5670;
            {7'd81,7'd71}:		p = 14'd5751;
            {7'd81,7'd72}:		p = 14'd5832;
            {7'd81,7'd73}:		p = 14'd5913;
            {7'd81,7'd74}:		p = 14'd5994;
            {7'd81,7'd75}:		p = 14'd6075;
            {7'd81,7'd76}:		p = 14'd6156;
            {7'd81,7'd77}:		p = 14'd6237;
            {7'd81,7'd78}:		p = 14'd6318;
            {7'd81,7'd79}:		p = 14'd6399;
            {7'd81,7'd80}:		p = 14'd6480;
            {7'd81,7'd81}:		p = 14'd6561;
            {7'd81,7'd82}:		p = 14'd6642;
            {7'd81,7'd83}:		p = 14'd6723;
            {7'd81,7'd84}:		p = 14'd6804;
            {7'd81,7'd85}:		p = 14'd6885;
            {7'd81,7'd86}:		p = 14'd6966;
            {7'd81,7'd87}:		p = 14'd7047;
            {7'd81,7'd88}:		p = 14'd7128;
            {7'd81,7'd89}:		p = 14'd7209;
            {7'd81,7'd90}:		p = 14'd7290;
            {7'd81,7'd91}:		p = 14'd7371;
            {7'd81,7'd92}:		p = 14'd7452;
            {7'd81,7'd93}:		p = 14'd7533;
            {7'd81,7'd94}:		p = 14'd7614;
            {7'd81,7'd95}:		p = 14'd7695;
            {7'd81,7'd96}:		p = 14'd7776;
            {7'd81,7'd97}:		p = 14'd7857;
            {7'd81,7'd98}:		p = 14'd7938;
            {7'd81,7'd99}:		p = 14'd8019;
            {7'd81,7'd100}:		p = 14'd8100;
            {7'd81,7'd101}:		p = 14'd8181;
            {7'd81,7'd102}:		p = 14'd8262;
            {7'd81,7'd103}:		p = 14'd8343;
            {7'd81,7'd104}:		p = 14'd8424;
            {7'd81,7'd105}:		p = 14'd8505;
            {7'd81,7'd106}:		p = 14'd8586;
            {7'd81,7'd107}:		p = 14'd8667;
            {7'd81,7'd108}:		p = 14'd8748;
            {7'd81,7'd109}:		p = 14'd8829;
            {7'd81,7'd110}:		p = 14'd8910;
            {7'd81,7'd111}:		p = 14'd8991;
            {7'd81,7'd112}:		p = 14'd9072;
            {7'd81,7'd113}:		p = 14'd9153;
            {7'd81,7'd114}:		p = 14'd9234;
            {7'd81,7'd115}:		p = 14'd9315;
            {7'd81,7'd116}:		p = 14'd9396;
            {7'd81,7'd117}:		p = 14'd9477;
            {7'd81,7'd118}:		p = 14'd9558;
            {7'd81,7'd119}:		p = 14'd9639;
            {7'd81,7'd120}:		p = 14'd9720;
            {7'd81,7'd121}:		p = 14'd9801;
            {7'd81,7'd122}:		p = 14'd9882;
            {7'd81,7'd123}:		p = 14'd9963;
            {7'd81,7'd124}:		p = 14'd10044;
            {7'd81,7'd125}:		p = 14'd10125;
            {7'd81,7'd126}:		p = 14'd10206;
            {7'd81,7'd127}:		p = 14'd10287;
            {7'd82,7'd0}:		p = 14'd0;
            {7'd82,7'd1}:		p = 14'd82;
            {7'd82,7'd2}:		p = 14'd164;
            {7'd82,7'd3}:		p = 14'd246;
            {7'd82,7'd4}:		p = 14'd328;
            {7'd82,7'd5}:		p = 14'd410;
            {7'd82,7'd6}:		p = 14'd492;
            {7'd82,7'd7}:		p = 14'd574;
            {7'd82,7'd8}:		p = 14'd656;
            {7'd82,7'd9}:		p = 14'd738;
            {7'd82,7'd10}:		p = 14'd820;
            {7'd82,7'd11}:		p = 14'd902;
            {7'd82,7'd12}:		p = 14'd984;
            {7'd82,7'd13}:		p = 14'd1066;
            {7'd82,7'd14}:		p = 14'd1148;
            {7'd82,7'd15}:		p = 14'd1230;
            {7'd82,7'd16}:		p = 14'd1312;
            {7'd82,7'd17}:		p = 14'd1394;
            {7'd82,7'd18}:		p = 14'd1476;
            {7'd82,7'd19}:		p = 14'd1558;
            {7'd82,7'd20}:		p = 14'd1640;
            {7'd82,7'd21}:		p = 14'd1722;
            {7'd82,7'd22}:		p = 14'd1804;
            {7'd82,7'd23}:		p = 14'd1886;
            {7'd82,7'd24}:		p = 14'd1968;
            {7'd82,7'd25}:		p = 14'd2050;
            {7'd82,7'd26}:		p = 14'd2132;
            {7'd82,7'd27}:		p = 14'd2214;
            {7'd82,7'd28}:		p = 14'd2296;
            {7'd82,7'd29}:		p = 14'd2378;
            {7'd82,7'd30}:		p = 14'd2460;
            {7'd82,7'd31}:		p = 14'd2542;
            {7'd82,7'd32}:		p = 14'd2624;
            {7'd82,7'd33}:		p = 14'd2706;
            {7'd82,7'd34}:		p = 14'd2788;
            {7'd82,7'd35}:		p = 14'd2870;
            {7'd82,7'd36}:		p = 14'd2952;
            {7'd82,7'd37}:		p = 14'd3034;
            {7'd82,7'd38}:		p = 14'd3116;
            {7'd82,7'd39}:		p = 14'd3198;
            {7'd82,7'd40}:		p = 14'd3280;
            {7'd82,7'd41}:		p = 14'd3362;
            {7'd82,7'd42}:		p = 14'd3444;
            {7'd82,7'd43}:		p = 14'd3526;
            {7'd82,7'd44}:		p = 14'd3608;
            {7'd82,7'd45}:		p = 14'd3690;
            {7'd82,7'd46}:		p = 14'd3772;
            {7'd82,7'd47}:		p = 14'd3854;
            {7'd82,7'd48}:		p = 14'd3936;
            {7'd82,7'd49}:		p = 14'd4018;
            {7'd82,7'd50}:		p = 14'd4100;
            {7'd82,7'd51}:		p = 14'd4182;
            {7'd82,7'd52}:		p = 14'd4264;
            {7'd82,7'd53}:		p = 14'd4346;
            {7'd82,7'd54}:		p = 14'd4428;
            {7'd82,7'd55}:		p = 14'd4510;
            {7'd82,7'd56}:		p = 14'd4592;
            {7'd82,7'd57}:		p = 14'd4674;
            {7'd82,7'd58}:		p = 14'd4756;
            {7'd82,7'd59}:		p = 14'd4838;
            {7'd82,7'd60}:		p = 14'd4920;
            {7'd82,7'd61}:		p = 14'd5002;
            {7'd82,7'd62}:		p = 14'd5084;
            {7'd82,7'd63}:		p = 14'd5166;
            {7'd82,7'd64}:		p = 14'd5248;
            {7'd82,7'd65}:		p = 14'd5330;
            {7'd82,7'd66}:		p = 14'd5412;
            {7'd82,7'd67}:		p = 14'd5494;
            {7'd82,7'd68}:		p = 14'd5576;
            {7'd82,7'd69}:		p = 14'd5658;
            {7'd82,7'd70}:		p = 14'd5740;
            {7'd82,7'd71}:		p = 14'd5822;
            {7'd82,7'd72}:		p = 14'd5904;
            {7'd82,7'd73}:		p = 14'd5986;
            {7'd82,7'd74}:		p = 14'd6068;
            {7'd82,7'd75}:		p = 14'd6150;
            {7'd82,7'd76}:		p = 14'd6232;
            {7'd82,7'd77}:		p = 14'd6314;
            {7'd82,7'd78}:		p = 14'd6396;
            {7'd82,7'd79}:		p = 14'd6478;
            {7'd82,7'd80}:		p = 14'd6560;
            {7'd82,7'd81}:		p = 14'd6642;
            {7'd82,7'd82}:		p = 14'd6724;
            {7'd82,7'd83}:		p = 14'd6806;
            {7'd82,7'd84}:		p = 14'd6888;
            {7'd82,7'd85}:		p = 14'd6970;
            {7'd82,7'd86}:		p = 14'd7052;
            {7'd82,7'd87}:		p = 14'd7134;
            {7'd82,7'd88}:		p = 14'd7216;
            {7'd82,7'd89}:		p = 14'd7298;
            {7'd82,7'd90}:		p = 14'd7380;
            {7'd82,7'd91}:		p = 14'd7462;
            {7'd82,7'd92}:		p = 14'd7544;
            {7'd82,7'd93}:		p = 14'd7626;
            {7'd82,7'd94}:		p = 14'd7708;
            {7'd82,7'd95}:		p = 14'd7790;
            {7'd82,7'd96}:		p = 14'd7872;
            {7'd82,7'd97}:		p = 14'd7954;
            {7'd82,7'd98}:		p = 14'd8036;
            {7'd82,7'd99}:		p = 14'd8118;
            {7'd82,7'd100}:		p = 14'd8200;
            {7'd82,7'd101}:		p = 14'd8282;
            {7'd82,7'd102}:		p = 14'd8364;
            {7'd82,7'd103}:		p = 14'd8446;
            {7'd82,7'd104}:		p = 14'd8528;
            {7'd82,7'd105}:		p = 14'd8610;
            {7'd82,7'd106}:		p = 14'd8692;
            {7'd82,7'd107}:		p = 14'd8774;
            {7'd82,7'd108}:		p = 14'd8856;
            {7'd82,7'd109}:		p = 14'd8938;
            {7'd82,7'd110}:		p = 14'd9020;
            {7'd82,7'd111}:		p = 14'd9102;
            {7'd82,7'd112}:		p = 14'd9184;
            {7'd82,7'd113}:		p = 14'd9266;
            {7'd82,7'd114}:		p = 14'd9348;
            {7'd82,7'd115}:		p = 14'd9430;
            {7'd82,7'd116}:		p = 14'd9512;
            {7'd82,7'd117}:		p = 14'd9594;
            {7'd82,7'd118}:		p = 14'd9676;
            {7'd82,7'd119}:		p = 14'd9758;
            {7'd82,7'd120}:		p = 14'd9840;
            {7'd82,7'd121}:		p = 14'd9922;
            {7'd82,7'd122}:		p = 14'd10004;
            {7'd82,7'd123}:		p = 14'd10086;
            {7'd82,7'd124}:		p = 14'd10168;
            {7'd82,7'd125}:		p = 14'd10250;
            {7'd82,7'd126}:		p = 14'd10332;
            {7'd82,7'd127}:		p = 14'd10414;
            {7'd83,7'd0}:		p = 14'd0;
            {7'd83,7'd1}:		p = 14'd83;
            {7'd83,7'd2}:		p = 14'd166;
            {7'd83,7'd3}:		p = 14'd249;
            {7'd83,7'd4}:		p = 14'd332;
            {7'd83,7'd5}:		p = 14'd415;
            {7'd83,7'd6}:		p = 14'd498;
            {7'd83,7'd7}:		p = 14'd581;
            {7'd83,7'd8}:		p = 14'd664;
            {7'd83,7'd9}:		p = 14'd747;
            {7'd83,7'd10}:		p = 14'd830;
            {7'd83,7'd11}:		p = 14'd913;
            {7'd83,7'd12}:		p = 14'd996;
            {7'd83,7'd13}:		p = 14'd1079;
            {7'd83,7'd14}:		p = 14'd1162;
            {7'd83,7'd15}:		p = 14'd1245;
            {7'd83,7'd16}:		p = 14'd1328;
            {7'd83,7'd17}:		p = 14'd1411;
            {7'd83,7'd18}:		p = 14'd1494;
            {7'd83,7'd19}:		p = 14'd1577;
            {7'd83,7'd20}:		p = 14'd1660;
            {7'd83,7'd21}:		p = 14'd1743;
            {7'd83,7'd22}:		p = 14'd1826;
            {7'd83,7'd23}:		p = 14'd1909;
            {7'd83,7'd24}:		p = 14'd1992;
            {7'd83,7'd25}:		p = 14'd2075;
            {7'd83,7'd26}:		p = 14'd2158;
            {7'd83,7'd27}:		p = 14'd2241;
            {7'd83,7'd28}:		p = 14'd2324;
            {7'd83,7'd29}:		p = 14'd2407;
            {7'd83,7'd30}:		p = 14'd2490;
            {7'd83,7'd31}:		p = 14'd2573;
            {7'd83,7'd32}:		p = 14'd2656;
            {7'd83,7'd33}:		p = 14'd2739;
            {7'd83,7'd34}:		p = 14'd2822;
            {7'd83,7'd35}:		p = 14'd2905;
            {7'd83,7'd36}:		p = 14'd2988;
            {7'd83,7'd37}:		p = 14'd3071;
            {7'd83,7'd38}:		p = 14'd3154;
            {7'd83,7'd39}:		p = 14'd3237;
            {7'd83,7'd40}:		p = 14'd3320;
            {7'd83,7'd41}:		p = 14'd3403;
            {7'd83,7'd42}:		p = 14'd3486;
            {7'd83,7'd43}:		p = 14'd3569;
            {7'd83,7'd44}:		p = 14'd3652;
            {7'd83,7'd45}:		p = 14'd3735;
            {7'd83,7'd46}:		p = 14'd3818;
            {7'd83,7'd47}:		p = 14'd3901;
            {7'd83,7'd48}:		p = 14'd3984;
            {7'd83,7'd49}:		p = 14'd4067;
            {7'd83,7'd50}:		p = 14'd4150;
            {7'd83,7'd51}:		p = 14'd4233;
            {7'd83,7'd52}:		p = 14'd4316;
            {7'd83,7'd53}:		p = 14'd4399;
            {7'd83,7'd54}:		p = 14'd4482;
            {7'd83,7'd55}:		p = 14'd4565;
            {7'd83,7'd56}:		p = 14'd4648;
            {7'd83,7'd57}:		p = 14'd4731;
            {7'd83,7'd58}:		p = 14'd4814;
            {7'd83,7'd59}:		p = 14'd4897;
            {7'd83,7'd60}:		p = 14'd4980;
            {7'd83,7'd61}:		p = 14'd5063;
            {7'd83,7'd62}:		p = 14'd5146;
            {7'd83,7'd63}:		p = 14'd5229;
            {7'd83,7'd64}:		p = 14'd5312;
            {7'd83,7'd65}:		p = 14'd5395;
            {7'd83,7'd66}:		p = 14'd5478;
            {7'd83,7'd67}:		p = 14'd5561;
            {7'd83,7'd68}:		p = 14'd5644;
            {7'd83,7'd69}:		p = 14'd5727;
            {7'd83,7'd70}:		p = 14'd5810;
            {7'd83,7'd71}:		p = 14'd5893;
            {7'd83,7'd72}:		p = 14'd5976;
            {7'd83,7'd73}:		p = 14'd6059;
            {7'd83,7'd74}:		p = 14'd6142;
            {7'd83,7'd75}:		p = 14'd6225;
            {7'd83,7'd76}:		p = 14'd6308;
            {7'd83,7'd77}:		p = 14'd6391;
            {7'd83,7'd78}:		p = 14'd6474;
            {7'd83,7'd79}:		p = 14'd6557;
            {7'd83,7'd80}:		p = 14'd6640;
            {7'd83,7'd81}:		p = 14'd6723;
            {7'd83,7'd82}:		p = 14'd6806;
            {7'd83,7'd83}:		p = 14'd6889;
            {7'd83,7'd84}:		p = 14'd6972;
            {7'd83,7'd85}:		p = 14'd7055;
            {7'd83,7'd86}:		p = 14'd7138;
            {7'd83,7'd87}:		p = 14'd7221;
            {7'd83,7'd88}:		p = 14'd7304;
            {7'd83,7'd89}:		p = 14'd7387;
            {7'd83,7'd90}:		p = 14'd7470;
            {7'd83,7'd91}:		p = 14'd7553;
            {7'd83,7'd92}:		p = 14'd7636;
            {7'd83,7'd93}:		p = 14'd7719;
            {7'd83,7'd94}:		p = 14'd7802;
            {7'd83,7'd95}:		p = 14'd7885;
            {7'd83,7'd96}:		p = 14'd7968;
            {7'd83,7'd97}:		p = 14'd8051;
            {7'd83,7'd98}:		p = 14'd8134;
            {7'd83,7'd99}:		p = 14'd8217;
            {7'd83,7'd100}:		p = 14'd8300;
            {7'd83,7'd101}:		p = 14'd8383;
            {7'd83,7'd102}:		p = 14'd8466;
            {7'd83,7'd103}:		p = 14'd8549;
            {7'd83,7'd104}:		p = 14'd8632;
            {7'd83,7'd105}:		p = 14'd8715;
            {7'd83,7'd106}:		p = 14'd8798;
            {7'd83,7'd107}:		p = 14'd8881;
            {7'd83,7'd108}:		p = 14'd8964;
            {7'd83,7'd109}:		p = 14'd9047;
            {7'd83,7'd110}:		p = 14'd9130;
            {7'd83,7'd111}:		p = 14'd9213;
            {7'd83,7'd112}:		p = 14'd9296;
            {7'd83,7'd113}:		p = 14'd9379;
            {7'd83,7'd114}:		p = 14'd9462;
            {7'd83,7'd115}:		p = 14'd9545;
            {7'd83,7'd116}:		p = 14'd9628;
            {7'd83,7'd117}:		p = 14'd9711;
            {7'd83,7'd118}:		p = 14'd9794;
            {7'd83,7'd119}:		p = 14'd9877;
            {7'd83,7'd120}:		p = 14'd9960;
            {7'd83,7'd121}:		p = 14'd10043;
            {7'd83,7'd122}:		p = 14'd10126;
            {7'd83,7'd123}:		p = 14'd10209;
            {7'd83,7'd124}:		p = 14'd10292;
            {7'd83,7'd125}:		p = 14'd10375;
            {7'd83,7'd126}:		p = 14'd10458;
            {7'd83,7'd127}:		p = 14'd10541;
            {7'd84,7'd0}:		p = 14'd0;
            {7'd84,7'd1}:		p = 14'd84;
            {7'd84,7'd2}:		p = 14'd168;
            {7'd84,7'd3}:		p = 14'd252;
            {7'd84,7'd4}:		p = 14'd336;
            {7'd84,7'd5}:		p = 14'd420;
            {7'd84,7'd6}:		p = 14'd504;
            {7'd84,7'd7}:		p = 14'd588;
            {7'd84,7'd8}:		p = 14'd672;
            {7'd84,7'd9}:		p = 14'd756;
            {7'd84,7'd10}:		p = 14'd840;
            {7'd84,7'd11}:		p = 14'd924;
            {7'd84,7'd12}:		p = 14'd1008;
            {7'd84,7'd13}:		p = 14'd1092;
            {7'd84,7'd14}:		p = 14'd1176;
            {7'd84,7'd15}:		p = 14'd1260;
            {7'd84,7'd16}:		p = 14'd1344;
            {7'd84,7'd17}:		p = 14'd1428;
            {7'd84,7'd18}:		p = 14'd1512;
            {7'd84,7'd19}:		p = 14'd1596;
            {7'd84,7'd20}:		p = 14'd1680;
            {7'd84,7'd21}:		p = 14'd1764;
            {7'd84,7'd22}:		p = 14'd1848;
            {7'd84,7'd23}:		p = 14'd1932;
            {7'd84,7'd24}:		p = 14'd2016;
            {7'd84,7'd25}:		p = 14'd2100;
            {7'd84,7'd26}:		p = 14'd2184;
            {7'd84,7'd27}:		p = 14'd2268;
            {7'd84,7'd28}:		p = 14'd2352;
            {7'd84,7'd29}:		p = 14'd2436;
            {7'd84,7'd30}:		p = 14'd2520;
            {7'd84,7'd31}:		p = 14'd2604;
            {7'd84,7'd32}:		p = 14'd2688;
            {7'd84,7'd33}:		p = 14'd2772;
            {7'd84,7'd34}:		p = 14'd2856;
            {7'd84,7'd35}:		p = 14'd2940;
            {7'd84,7'd36}:		p = 14'd3024;
            {7'd84,7'd37}:		p = 14'd3108;
            {7'd84,7'd38}:		p = 14'd3192;
            {7'd84,7'd39}:		p = 14'd3276;
            {7'd84,7'd40}:		p = 14'd3360;
            {7'd84,7'd41}:		p = 14'd3444;
            {7'd84,7'd42}:		p = 14'd3528;
            {7'd84,7'd43}:		p = 14'd3612;
            {7'd84,7'd44}:		p = 14'd3696;
            {7'd84,7'd45}:		p = 14'd3780;
            {7'd84,7'd46}:		p = 14'd3864;
            {7'd84,7'd47}:		p = 14'd3948;
            {7'd84,7'd48}:		p = 14'd4032;
            {7'd84,7'd49}:		p = 14'd4116;
            {7'd84,7'd50}:		p = 14'd4200;
            {7'd84,7'd51}:		p = 14'd4284;
            {7'd84,7'd52}:		p = 14'd4368;
            {7'd84,7'd53}:		p = 14'd4452;
            {7'd84,7'd54}:		p = 14'd4536;
            {7'd84,7'd55}:		p = 14'd4620;
            {7'd84,7'd56}:		p = 14'd4704;
            {7'd84,7'd57}:		p = 14'd4788;
            {7'd84,7'd58}:		p = 14'd4872;
            {7'd84,7'd59}:		p = 14'd4956;
            {7'd84,7'd60}:		p = 14'd5040;
            {7'd84,7'd61}:		p = 14'd5124;
            {7'd84,7'd62}:		p = 14'd5208;
            {7'd84,7'd63}:		p = 14'd5292;
            {7'd84,7'd64}:		p = 14'd5376;
            {7'd84,7'd65}:		p = 14'd5460;
            {7'd84,7'd66}:		p = 14'd5544;
            {7'd84,7'd67}:		p = 14'd5628;
            {7'd84,7'd68}:		p = 14'd5712;
            {7'd84,7'd69}:		p = 14'd5796;
            {7'd84,7'd70}:		p = 14'd5880;
            {7'd84,7'd71}:		p = 14'd5964;
            {7'd84,7'd72}:		p = 14'd6048;
            {7'd84,7'd73}:		p = 14'd6132;
            {7'd84,7'd74}:		p = 14'd6216;
            {7'd84,7'd75}:		p = 14'd6300;
            {7'd84,7'd76}:		p = 14'd6384;
            {7'd84,7'd77}:		p = 14'd6468;
            {7'd84,7'd78}:		p = 14'd6552;
            {7'd84,7'd79}:		p = 14'd6636;
            {7'd84,7'd80}:		p = 14'd6720;
            {7'd84,7'd81}:		p = 14'd6804;
            {7'd84,7'd82}:		p = 14'd6888;
            {7'd84,7'd83}:		p = 14'd6972;
            {7'd84,7'd84}:		p = 14'd7056;
            {7'd84,7'd85}:		p = 14'd7140;
            {7'd84,7'd86}:		p = 14'd7224;
            {7'd84,7'd87}:		p = 14'd7308;
            {7'd84,7'd88}:		p = 14'd7392;
            {7'd84,7'd89}:		p = 14'd7476;
            {7'd84,7'd90}:		p = 14'd7560;
            {7'd84,7'd91}:		p = 14'd7644;
            {7'd84,7'd92}:		p = 14'd7728;
            {7'd84,7'd93}:		p = 14'd7812;
            {7'd84,7'd94}:		p = 14'd7896;
            {7'd84,7'd95}:		p = 14'd7980;
            {7'd84,7'd96}:		p = 14'd8064;
            {7'd84,7'd97}:		p = 14'd8148;
            {7'd84,7'd98}:		p = 14'd8232;
            {7'd84,7'd99}:		p = 14'd8316;
            {7'd84,7'd100}:		p = 14'd8400;
            {7'd84,7'd101}:		p = 14'd8484;
            {7'd84,7'd102}:		p = 14'd8568;
            {7'd84,7'd103}:		p = 14'd8652;
            {7'd84,7'd104}:		p = 14'd8736;
            {7'd84,7'd105}:		p = 14'd8820;
            {7'd84,7'd106}:		p = 14'd8904;
            {7'd84,7'd107}:		p = 14'd8988;
            {7'd84,7'd108}:		p = 14'd9072;
            {7'd84,7'd109}:		p = 14'd9156;
            {7'd84,7'd110}:		p = 14'd9240;
            {7'd84,7'd111}:		p = 14'd9324;
            {7'd84,7'd112}:		p = 14'd9408;
            {7'd84,7'd113}:		p = 14'd9492;
            {7'd84,7'd114}:		p = 14'd9576;
            {7'd84,7'd115}:		p = 14'd9660;
            {7'd84,7'd116}:		p = 14'd9744;
            {7'd84,7'd117}:		p = 14'd9828;
            {7'd84,7'd118}:		p = 14'd9912;
            {7'd84,7'd119}:		p = 14'd9996;
            {7'd84,7'd120}:		p = 14'd10080;
            {7'd84,7'd121}:		p = 14'd10164;
            {7'd84,7'd122}:		p = 14'd10248;
            {7'd84,7'd123}:		p = 14'd10332;
            {7'd84,7'd124}:		p = 14'd10416;
            {7'd84,7'd125}:		p = 14'd10500;
            {7'd84,7'd126}:		p = 14'd10584;
            {7'd84,7'd127}:		p = 14'd10668;
            {7'd85,7'd0}:		p = 14'd0;
            {7'd85,7'd1}:		p = 14'd85;
            {7'd85,7'd2}:		p = 14'd170;
            {7'd85,7'd3}:		p = 14'd255;
            {7'd85,7'd4}:		p = 14'd340;
            {7'd85,7'd5}:		p = 14'd425;
            {7'd85,7'd6}:		p = 14'd510;
            {7'd85,7'd7}:		p = 14'd595;
            {7'd85,7'd8}:		p = 14'd680;
            {7'd85,7'd9}:		p = 14'd765;
            {7'd85,7'd10}:		p = 14'd850;
            {7'd85,7'd11}:		p = 14'd935;
            {7'd85,7'd12}:		p = 14'd1020;
            {7'd85,7'd13}:		p = 14'd1105;
            {7'd85,7'd14}:		p = 14'd1190;
            {7'd85,7'd15}:		p = 14'd1275;
            {7'd85,7'd16}:		p = 14'd1360;
            {7'd85,7'd17}:		p = 14'd1445;
            {7'd85,7'd18}:		p = 14'd1530;
            {7'd85,7'd19}:		p = 14'd1615;
            {7'd85,7'd20}:		p = 14'd1700;
            {7'd85,7'd21}:		p = 14'd1785;
            {7'd85,7'd22}:		p = 14'd1870;
            {7'd85,7'd23}:		p = 14'd1955;
            {7'd85,7'd24}:		p = 14'd2040;
            {7'd85,7'd25}:		p = 14'd2125;
            {7'd85,7'd26}:		p = 14'd2210;
            {7'd85,7'd27}:		p = 14'd2295;
            {7'd85,7'd28}:		p = 14'd2380;
            {7'd85,7'd29}:		p = 14'd2465;
            {7'd85,7'd30}:		p = 14'd2550;
            {7'd85,7'd31}:		p = 14'd2635;
            {7'd85,7'd32}:		p = 14'd2720;
            {7'd85,7'd33}:		p = 14'd2805;
            {7'd85,7'd34}:		p = 14'd2890;
            {7'd85,7'd35}:		p = 14'd2975;
            {7'd85,7'd36}:		p = 14'd3060;
            {7'd85,7'd37}:		p = 14'd3145;
            {7'd85,7'd38}:		p = 14'd3230;
            {7'd85,7'd39}:		p = 14'd3315;
            {7'd85,7'd40}:		p = 14'd3400;
            {7'd85,7'd41}:		p = 14'd3485;
            {7'd85,7'd42}:		p = 14'd3570;
            {7'd85,7'd43}:		p = 14'd3655;
            {7'd85,7'd44}:		p = 14'd3740;
            {7'd85,7'd45}:		p = 14'd3825;
            {7'd85,7'd46}:		p = 14'd3910;
            {7'd85,7'd47}:		p = 14'd3995;
            {7'd85,7'd48}:		p = 14'd4080;
            {7'd85,7'd49}:		p = 14'd4165;
            {7'd85,7'd50}:		p = 14'd4250;
            {7'd85,7'd51}:		p = 14'd4335;
            {7'd85,7'd52}:		p = 14'd4420;
            {7'd85,7'd53}:		p = 14'd4505;
            {7'd85,7'd54}:		p = 14'd4590;
            {7'd85,7'd55}:		p = 14'd4675;
            {7'd85,7'd56}:		p = 14'd4760;
            {7'd85,7'd57}:		p = 14'd4845;
            {7'd85,7'd58}:		p = 14'd4930;
            {7'd85,7'd59}:		p = 14'd5015;
            {7'd85,7'd60}:		p = 14'd5100;
            {7'd85,7'd61}:		p = 14'd5185;
            {7'd85,7'd62}:		p = 14'd5270;
            {7'd85,7'd63}:		p = 14'd5355;
            {7'd85,7'd64}:		p = 14'd5440;
            {7'd85,7'd65}:		p = 14'd5525;
            {7'd85,7'd66}:		p = 14'd5610;
            {7'd85,7'd67}:		p = 14'd5695;
            {7'd85,7'd68}:		p = 14'd5780;
            {7'd85,7'd69}:		p = 14'd5865;
            {7'd85,7'd70}:		p = 14'd5950;
            {7'd85,7'd71}:		p = 14'd6035;
            {7'd85,7'd72}:		p = 14'd6120;
            {7'd85,7'd73}:		p = 14'd6205;
            {7'd85,7'd74}:		p = 14'd6290;
            {7'd85,7'd75}:		p = 14'd6375;
            {7'd85,7'd76}:		p = 14'd6460;
            {7'd85,7'd77}:		p = 14'd6545;
            {7'd85,7'd78}:		p = 14'd6630;
            {7'd85,7'd79}:		p = 14'd6715;
            {7'd85,7'd80}:		p = 14'd6800;
            {7'd85,7'd81}:		p = 14'd6885;
            {7'd85,7'd82}:		p = 14'd6970;
            {7'd85,7'd83}:		p = 14'd7055;
            {7'd85,7'd84}:		p = 14'd7140;
            {7'd85,7'd85}:		p = 14'd7225;
            {7'd85,7'd86}:		p = 14'd7310;
            {7'd85,7'd87}:		p = 14'd7395;
            {7'd85,7'd88}:		p = 14'd7480;
            {7'd85,7'd89}:		p = 14'd7565;
            {7'd85,7'd90}:		p = 14'd7650;
            {7'd85,7'd91}:		p = 14'd7735;
            {7'd85,7'd92}:		p = 14'd7820;
            {7'd85,7'd93}:		p = 14'd7905;
            {7'd85,7'd94}:		p = 14'd7990;
            {7'd85,7'd95}:		p = 14'd8075;
            {7'd85,7'd96}:		p = 14'd8160;
            {7'd85,7'd97}:		p = 14'd8245;
            {7'd85,7'd98}:		p = 14'd8330;
            {7'd85,7'd99}:		p = 14'd8415;
            {7'd85,7'd100}:		p = 14'd8500;
            {7'd85,7'd101}:		p = 14'd8585;
            {7'd85,7'd102}:		p = 14'd8670;
            {7'd85,7'd103}:		p = 14'd8755;
            {7'd85,7'd104}:		p = 14'd8840;
            {7'd85,7'd105}:		p = 14'd8925;
            {7'd85,7'd106}:		p = 14'd9010;
            {7'd85,7'd107}:		p = 14'd9095;
            {7'd85,7'd108}:		p = 14'd9180;
            {7'd85,7'd109}:		p = 14'd9265;
            {7'd85,7'd110}:		p = 14'd9350;
            {7'd85,7'd111}:		p = 14'd9435;
            {7'd85,7'd112}:		p = 14'd9520;
            {7'd85,7'd113}:		p = 14'd9605;
            {7'd85,7'd114}:		p = 14'd9690;
            {7'd85,7'd115}:		p = 14'd9775;
            {7'd85,7'd116}:		p = 14'd9860;
            {7'd85,7'd117}:		p = 14'd9945;
            {7'd85,7'd118}:		p = 14'd10030;
            {7'd85,7'd119}:		p = 14'd10115;
            {7'd85,7'd120}:		p = 14'd10200;
            {7'd85,7'd121}:		p = 14'd10285;
            {7'd85,7'd122}:		p = 14'd10370;
            {7'd85,7'd123}:		p = 14'd10455;
            {7'd85,7'd124}:		p = 14'd10540;
            {7'd85,7'd125}:		p = 14'd10625;
            {7'd85,7'd126}:		p = 14'd10710;
            {7'd85,7'd127}:		p = 14'd10795;
            {7'd86,7'd0}:		p = 14'd0;
            {7'd86,7'd1}:		p = 14'd86;
            {7'd86,7'd2}:		p = 14'd172;
            {7'd86,7'd3}:		p = 14'd258;
            {7'd86,7'd4}:		p = 14'd344;
            {7'd86,7'd5}:		p = 14'd430;
            {7'd86,7'd6}:		p = 14'd516;
            {7'd86,7'd7}:		p = 14'd602;
            {7'd86,7'd8}:		p = 14'd688;
            {7'd86,7'd9}:		p = 14'd774;
            {7'd86,7'd10}:		p = 14'd860;
            {7'd86,7'd11}:		p = 14'd946;
            {7'd86,7'd12}:		p = 14'd1032;
            {7'd86,7'd13}:		p = 14'd1118;
            {7'd86,7'd14}:		p = 14'd1204;
            {7'd86,7'd15}:		p = 14'd1290;
            {7'd86,7'd16}:		p = 14'd1376;
            {7'd86,7'd17}:		p = 14'd1462;
            {7'd86,7'd18}:		p = 14'd1548;
            {7'd86,7'd19}:		p = 14'd1634;
            {7'd86,7'd20}:		p = 14'd1720;
            {7'd86,7'd21}:		p = 14'd1806;
            {7'd86,7'd22}:		p = 14'd1892;
            {7'd86,7'd23}:		p = 14'd1978;
            {7'd86,7'd24}:		p = 14'd2064;
            {7'd86,7'd25}:		p = 14'd2150;
            {7'd86,7'd26}:		p = 14'd2236;
            {7'd86,7'd27}:		p = 14'd2322;
            {7'd86,7'd28}:		p = 14'd2408;
            {7'd86,7'd29}:		p = 14'd2494;
            {7'd86,7'd30}:		p = 14'd2580;
            {7'd86,7'd31}:		p = 14'd2666;
            {7'd86,7'd32}:		p = 14'd2752;
            {7'd86,7'd33}:		p = 14'd2838;
            {7'd86,7'd34}:		p = 14'd2924;
            {7'd86,7'd35}:		p = 14'd3010;
            {7'd86,7'd36}:		p = 14'd3096;
            {7'd86,7'd37}:		p = 14'd3182;
            {7'd86,7'd38}:		p = 14'd3268;
            {7'd86,7'd39}:		p = 14'd3354;
            {7'd86,7'd40}:		p = 14'd3440;
            {7'd86,7'd41}:		p = 14'd3526;
            {7'd86,7'd42}:		p = 14'd3612;
            {7'd86,7'd43}:		p = 14'd3698;
            {7'd86,7'd44}:		p = 14'd3784;
            {7'd86,7'd45}:		p = 14'd3870;
            {7'd86,7'd46}:		p = 14'd3956;
            {7'd86,7'd47}:		p = 14'd4042;
            {7'd86,7'd48}:		p = 14'd4128;
            {7'd86,7'd49}:		p = 14'd4214;
            {7'd86,7'd50}:		p = 14'd4300;
            {7'd86,7'd51}:		p = 14'd4386;
            {7'd86,7'd52}:		p = 14'd4472;
            {7'd86,7'd53}:		p = 14'd4558;
            {7'd86,7'd54}:		p = 14'd4644;
            {7'd86,7'd55}:		p = 14'd4730;
            {7'd86,7'd56}:		p = 14'd4816;
            {7'd86,7'd57}:		p = 14'd4902;
            {7'd86,7'd58}:		p = 14'd4988;
            {7'd86,7'd59}:		p = 14'd5074;
            {7'd86,7'd60}:		p = 14'd5160;
            {7'd86,7'd61}:		p = 14'd5246;
            {7'd86,7'd62}:		p = 14'd5332;
            {7'd86,7'd63}:		p = 14'd5418;
            {7'd86,7'd64}:		p = 14'd5504;
            {7'd86,7'd65}:		p = 14'd5590;
            {7'd86,7'd66}:		p = 14'd5676;
            {7'd86,7'd67}:		p = 14'd5762;
            {7'd86,7'd68}:		p = 14'd5848;
            {7'd86,7'd69}:		p = 14'd5934;
            {7'd86,7'd70}:		p = 14'd6020;
            {7'd86,7'd71}:		p = 14'd6106;
            {7'd86,7'd72}:		p = 14'd6192;
            {7'd86,7'd73}:		p = 14'd6278;
            {7'd86,7'd74}:		p = 14'd6364;
            {7'd86,7'd75}:		p = 14'd6450;
            {7'd86,7'd76}:		p = 14'd6536;
            {7'd86,7'd77}:		p = 14'd6622;
            {7'd86,7'd78}:		p = 14'd6708;
            {7'd86,7'd79}:		p = 14'd6794;
            {7'd86,7'd80}:		p = 14'd6880;
            {7'd86,7'd81}:		p = 14'd6966;
            {7'd86,7'd82}:		p = 14'd7052;
            {7'd86,7'd83}:		p = 14'd7138;
            {7'd86,7'd84}:		p = 14'd7224;
            {7'd86,7'd85}:		p = 14'd7310;
            {7'd86,7'd86}:		p = 14'd7396;
            {7'd86,7'd87}:		p = 14'd7482;
            {7'd86,7'd88}:		p = 14'd7568;
            {7'd86,7'd89}:		p = 14'd7654;
            {7'd86,7'd90}:		p = 14'd7740;
            {7'd86,7'd91}:		p = 14'd7826;
            {7'd86,7'd92}:		p = 14'd7912;
            {7'd86,7'd93}:		p = 14'd7998;
            {7'd86,7'd94}:		p = 14'd8084;
            {7'd86,7'd95}:		p = 14'd8170;
            {7'd86,7'd96}:		p = 14'd8256;
            {7'd86,7'd97}:		p = 14'd8342;
            {7'd86,7'd98}:		p = 14'd8428;
            {7'd86,7'd99}:		p = 14'd8514;
            {7'd86,7'd100}:		p = 14'd8600;
            {7'd86,7'd101}:		p = 14'd8686;
            {7'd86,7'd102}:		p = 14'd8772;
            {7'd86,7'd103}:		p = 14'd8858;
            {7'd86,7'd104}:		p = 14'd8944;
            {7'd86,7'd105}:		p = 14'd9030;
            {7'd86,7'd106}:		p = 14'd9116;
            {7'd86,7'd107}:		p = 14'd9202;
            {7'd86,7'd108}:		p = 14'd9288;
            {7'd86,7'd109}:		p = 14'd9374;
            {7'd86,7'd110}:		p = 14'd9460;
            {7'd86,7'd111}:		p = 14'd9546;
            {7'd86,7'd112}:		p = 14'd9632;
            {7'd86,7'd113}:		p = 14'd9718;
            {7'd86,7'd114}:		p = 14'd9804;
            {7'd86,7'd115}:		p = 14'd9890;
            {7'd86,7'd116}:		p = 14'd9976;
            {7'd86,7'd117}:		p = 14'd10062;
            {7'd86,7'd118}:		p = 14'd10148;
            {7'd86,7'd119}:		p = 14'd10234;
            {7'd86,7'd120}:		p = 14'd10320;
            {7'd86,7'd121}:		p = 14'd10406;
            {7'd86,7'd122}:		p = 14'd10492;
            {7'd86,7'd123}:		p = 14'd10578;
            {7'd86,7'd124}:		p = 14'd10664;
            {7'd86,7'd125}:		p = 14'd10750;
            {7'd86,7'd126}:		p = 14'd10836;
            {7'd86,7'd127}:		p = 14'd10922;
            {7'd87,7'd0}:		p = 14'd0;
            {7'd87,7'd1}:		p = 14'd87;
            {7'd87,7'd2}:		p = 14'd174;
            {7'd87,7'd3}:		p = 14'd261;
            {7'd87,7'd4}:		p = 14'd348;
            {7'd87,7'd5}:		p = 14'd435;
            {7'd87,7'd6}:		p = 14'd522;
            {7'd87,7'd7}:		p = 14'd609;
            {7'd87,7'd8}:		p = 14'd696;
            {7'd87,7'd9}:		p = 14'd783;
            {7'd87,7'd10}:		p = 14'd870;
            {7'd87,7'd11}:		p = 14'd957;
            {7'd87,7'd12}:		p = 14'd1044;
            {7'd87,7'd13}:		p = 14'd1131;
            {7'd87,7'd14}:		p = 14'd1218;
            {7'd87,7'd15}:		p = 14'd1305;
            {7'd87,7'd16}:		p = 14'd1392;
            {7'd87,7'd17}:		p = 14'd1479;
            {7'd87,7'd18}:		p = 14'd1566;
            {7'd87,7'd19}:		p = 14'd1653;
            {7'd87,7'd20}:		p = 14'd1740;
            {7'd87,7'd21}:		p = 14'd1827;
            {7'd87,7'd22}:		p = 14'd1914;
            {7'd87,7'd23}:		p = 14'd2001;
            {7'd87,7'd24}:		p = 14'd2088;
            {7'd87,7'd25}:		p = 14'd2175;
            {7'd87,7'd26}:		p = 14'd2262;
            {7'd87,7'd27}:		p = 14'd2349;
            {7'd87,7'd28}:		p = 14'd2436;
            {7'd87,7'd29}:		p = 14'd2523;
            {7'd87,7'd30}:		p = 14'd2610;
            {7'd87,7'd31}:		p = 14'd2697;
            {7'd87,7'd32}:		p = 14'd2784;
            {7'd87,7'd33}:		p = 14'd2871;
            {7'd87,7'd34}:		p = 14'd2958;
            {7'd87,7'd35}:		p = 14'd3045;
            {7'd87,7'd36}:		p = 14'd3132;
            {7'd87,7'd37}:		p = 14'd3219;
            {7'd87,7'd38}:		p = 14'd3306;
            {7'd87,7'd39}:		p = 14'd3393;
            {7'd87,7'd40}:		p = 14'd3480;
            {7'd87,7'd41}:		p = 14'd3567;
            {7'd87,7'd42}:		p = 14'd3654;
            {7'd87,7'd43}:		p = 14'd3741;
            {7'd87,7'd44}:		p = 14'd3828;
            {7'd87,7'd45}:		p = 14'd3915;
            {7'd87,7'd46}:		p = 14'd4002;
            {7'd87,7'd47}:		p = 14'd4089;
            {7'd87,7'd48}:		p = 14'd4176;
            {7'd87,7'd49}:		p = 14'd4263;
            {7'd87,7'd50}:		p = 14'd4350;
            {7'd87,7'd51}:		p = 14'd4437;
            {7'd87,7'd52}:		p = 14'd4524;
            {7'd87,7'd53}:		p = 14'd4611;
            {7'd87,7'd54}:		p = 14'd4698;
            {7'd87,7'd55}:		p = 14'd4785;
            {7'd87,7'd56}:		p = 14'd4872;
            {7'd87,7'd57}:		p = 14'd4959;
            {7'd87,7'd58}:		p = 14'd5046;
            {7'd87,7'd59}:		p = 14'd5133;
            {7'd87,7'd60}:		p = 14'd5220;
            {7'd87,7'd61}:		p = 14'd5307;
            {7'd87,7'd62}:		p = 14'd5394;
            {7'd87,7'd63}:		p = 14'd5481;
            {7'd87,7'd64}:		p = 14'd5568;
            {7'd87,7'd65}:		p = 14'd5655;
            {7'd87,7'd66}:		p = 14'd5742;
            {7'd87,7'd67}:		p = 14'd5829;
            {7'd87,7'd68}:		p = 14'd5916;
            {7'd87,7'd69}:		p = 14'd6003;
            {7'd87,7'd70}:		p = 14'd6090;
            {7'd87,7'd71}:		p = 14'd6177;
            {7'd87,7'd72}:		p = 14'd6264;
            {7'd87,7'd73}:		p = 14'd6351;
            {7'd87,7'd74}:		p = 14'd6438;
            {7'd87,7'd75}:		p = 14'd6525;
            {7'd87,7'd76}:		p = 14'd6612;
            {7'd87,7'd77}:		p = 14'd6699;
            {7'd87,7'd78}:		p = 14'd6786;
            {7'd87,7'd79}:		p = 14'd6873;
            {7'd87,7'd80}:		p = 14'd6960;
            {7'd87,7'd81}:		p = 14'd7047;
            {7'd87,7'd82}:		p = 14'd7134;
            {7'd87,7'd83}:		p = 14'd7221;
            {7'd87,7'd84}:		p = 14'd7308;
            {7'd87,7'd85}:		p = 14'd7395;
            {7'd87,7'd86}:		p = 14'd7482;
            {7'd87,7'd87}:		p = 14'd7569;
            {7'd87,7'd88}:		p = 14'd7656;
            {7'd87,7'd89}:		p = 14'd7743;
            {7'd87,7'd90}:		p = 14'd7830;
            {7'd87,7'd91}:		p = 14'd7917;
            {7'd87,7'd92}:		p = 14'd8004;
            {7'd87,7'd93}:		p = 14'd8091;
            {7'd87,7'd94}:		p = 14'd8178;
            {7'd87,7'd95}:		p = 14'd8265;
            {7'd87,7'd96}:		p = 14'd8352;
            {7'd87,7'd97}:		p = 14'd8439;
            {7'd87,7'd98}:		p = 14'd8526;
            {7'd87,7'd99}:		p = 14'd8613;
            {7'd87,7'd100}:		p = 14'd8700;
            {7'd87,7'd101}:		p = 14'd8787;
            {7'd87,7'd102}:		p = 14'd8874;
            {7'd87,7'd103}:		p = 14'd8961;
            {7'd87,7'd104}:		p = 14'd9048;
            {7'd87,7'd105}:		p = 14'd9135;
            {7'd87,7'd106}:		p = 14'd9222;
            {7'd87,7'd107}:		p = 14'd9309;
            {7'd87,7'd108}:		p = 14'd9396;
            {7'd87,7'd109}:		p = 14'd9483;
            {7'd87,7'd110}:		p = 14'd9570;
            {7'd87,7'd111}:		p = 14'd9657;
            {7'd87,7'd112}:		p = 14'd9744;
            {7'd87,7'd113}:		p = 14'd9831;
            {7'd87,7'd114}:		p = 14'd9918;
            {7'd87,7'd115}:		p = 14'd10005;
            {7'd87,7'd116}:		p = 14'd10092;
            {7'd87,7'd117}:		p = 14'd10179;
            {7'd87,7'd118}:		p = 14'd10266;
            {7'd87,7'd119}:		p = 14'd10353;
            {7'd87,7'd120}:		p = 14'd10440;
            {7'd87,7'd121}:		p = 14'd10527;
            {7'd87,7'd122}:		p = 14'd10614;
            {7'd87,7'd123}:		p = 14'd10701;
            {7'd87,7'd124}:		p = 14'd10788;
            {7'd87,7'd125}:		p = 14'd10875;
            {7'd87,7'd126}:		p = 14'd10962;
            {7'd87,7'd127}:		p = 14'd11049;
            {7'd88,7'd0}:		p = 14'd0;
            {7'd88,7'd1}:		p = 14'd88;
            {7'd88,7'd2}:		p = 14'd176;
            {7'd88,7'd3}:		p = 14'd264;
            {7'd88,7'd4}:		p = 14'd352;
            {7'd88,7'd5}:		p = 14'd440;
            {7'd88,7'd6}:		p = 14'd528;
            {7'd88,7'd7}:		p = 14'd616;
            {7'd88,7'd8}:		p = 14'd704;
            {7'd88,7'd9}:		p = 14'd792;
            {7'd88,7'd10}:		p = 14'd880;
            {7'd88,7'd11}:		p = 14'd968;
            {7'd88,7'd12}:		p = 14'd1056;
            {7'd88,7'd13}:		p = 14'd1144;
            {7'd88,7'd14}:		p = 14'd1232;
            {7'd88,7'd15}:		p = 14'd1320;
            {7'd88,7'd16}:		p = 14'd1408;
            {7'd88,7'd17}:		p = 14'd1496;
            {7'd88,7'd18}:		p = 14'd1584;
            {7'd88,7'd19}:		p = 14'd1672;
            {7'd88,7'd20}:		p = 14'd1760;
            {7'd88,7'd21}:		p = 14'd1848;
            {7'd88,7'd22}:		p = 14'd1936;
            {7'd88,7'd23}:		p = 14'd2024;
            {7'd88,7'd24}:		p = 14'd2112;
            {7'd88,7'd25}:		p = 14'd2200;
            {7'd88,7'd26}:		p = 14'd2288;
            {7'd88,7'd27}:		p = 14'd2376;
            {7'd88,7'd28}:		p = 14'd2464;
            {7'd88,7'd29}:		p = 14'd2552;
            {7'd88,7'd30}:		p = 14'd2640;
            {7'd88,7'd31}:		p = 14'd2728;
            {7'd88,7'd32}:		p = 14'd2816;
            {7'd88,7'd33}:		p = 14'd2904;
            {7'd88,7'd34}:		p = 14'd2992;
            {7'd88,7'd35}:		p = 14'd3080;
            {7'd88,7'd36}:		p = 14'd3168;
            {7'd88,7'd37}:		p = 14'd3256;
            {7'd88,7'd38}:		p = 14'd3344;
            {7'd88,7'd39}:		p = 14'd3432;
            {7'd88,7'd40}:		p = 14'd3520;
            {7'd88,7'd41}:		p = 14'd3608;
            {7'd88,7'd42}:		p = 14'd3696;
            {7'd88,7'd43}:		p = 14'd3784;
            {7'd88,7'd44}:		p = 14'd3872;
            {7'd88,7'd45}:		p = 14'd3960;
            {7'd88,7'd46}:		p = 14'd4048;
            {7'd88,7'd47}:		p = 14'd4136;
            {7'd88,7'd48}:		p = 14'd4224;
            {7'd88,7'd49}:		p = 14'd4312;
            {7'd88,7'd50}:		p = 14'd4400;
            {7'd88,7'd51}:		p = 14'd4488;
            {7'd88,7'd52}:		p = 14'd4576;
            {7'd88,7'd53}:		p = 14'd4664;
            {7'd88,7'd54}:		p = 14'd4752;
            {7'd88,7'd55}:		p = 14'd4840;
            {7'd88,7'd56}:		p = 14'd4928;
            {7'd88,7'd57}:		p = 14'd5016;
            {7'd88,7'd58}:		p = 14'd5104;
            {7'd88,7'd59}:		p = 14'd5192;
            {7'd88,7'd60}:		p = 14'd5280;
            {7'd88,7'd61}:		p = 14'd5368;
            {7'd88,7'd62}:		p = 14'd5456;
            {7'd88,7'd63}:		p = 14'd5544;
            {7'd88,7'd64}:		p = 14'd5632;
            {7'd88,7'd65}:		p = 14'd5720;
            {7'd88,7'd66}:		p = 14'd5808;
            {7'd88,7'd67}:		p = 14'd5896;
            {7'd88,7'd68}:		p = 14'd5984;
            {7'd88,7'd69}:		p = 14'd6072;
            {7'd88,7'd70}:		p = 14'd6160;
            {7'd88,7'd71}:		p = 14'd6248;
            {7'd88,7'd72}:		p = 14'd6336;
            {7'd88,7'd73}:		p = 14'd6424;
            {7'd88,7'd74}:		p = 14'd6512;
            {7'd88,7'd75}:		p = 14'd6600;
            {7'd88,7'd76}:		p = 14'd6688;
            {7'd88,7'd77}:		p = 14'd6776;
            {7'd88,7'd78}:		p = 14'd6864;
            {7'd88,7'd79}:		p = 14'd6952;
            {7'd88,7'd80}:		p = 14'd7040;
            {7'd88,7'd81}:		p = 14'd7128;
            {7'd88,7'd82}:		p = 14'd7216;
            {7'd88,7'd83}:		p = 14'd7304;
            {7'd88,7'd84}:		p = 14'd7392;
            {7'd88,7'd85}:		p = 14'd7480;
            {7'd88,7'd86}:		p = 14'd7568;
            {7'd88,7'd87}:		p = 14'd7656;
            {7'd88,7'd88}:		p = 14'd7744;
            {7'd88,7'd89}:		p = 14'd7832;
            {7'd88,7'd90}:		p = 14'd7920;
            {7'd88,7'd91}:		p = 14'd8008;
            {7'd88,7'd92}:		p = 14'd8096;
            {7'd88,7'd93}:		p = 14'd8184;
            {7'd88,7'd94}:		p = 14'd8272;
            {7'd88,7'd95}:		p = 14'd8360;
            {7'd88,7'd96}:		p = 14'd8448;
            {7'd88,7'd97}:		p = 14'd8536;
            {7'd88,7'd98}:		p = 14'd8624;
            {7'd88,7'd99}:		p = 14'd8712;
            {7'd88,7'd100}:		p = 14'd8800;
            {7'd88,7'd101}:		p = 14'd8888;
            {7'd88,7'd102}:		p = 14'd8976;
            {7'd88,7'd103}:		p = 14'd9064;
            {7'd88,7'd104}:		p = 14'd9152;
            {7'd88,7'd105}:		p = 14'd9240;
            {7'd88,7'd106}:		p = 14'd9328;
            {7'd88,7'd107}:		p = 14'd9416;
            {7'd88,7'd108}:		p = 14'd9504;
            {7'd88,7'd109}:		p = 14'd9592;
            {7'd88,7'd110}:		p = 14'd9680;
            {7'd88,7'd111}:		p = 14'd9768;
            {7'd88,7'd112}:		p = 14'd9856;
            {7'd88,7'd113}:		p = 14'd9944;
            {7'd88,7'd114}:		p = 14'd10032;
            {7'd88,7'd115}:		p = 14'd10120;
            {7'd88,7'd116}:		p = 14'd10208;
            {7'd88,7'd117}:		p = 14'd10296;
            {7'd88,7'd118}:		p = 14'd10384;
            {7'd88,7'd119}:		p = 14'd10472;
            {7'd88,7'd120}:		p = 14'd10560;
            {7'd88,7'd121}:		p = 14'd10648;
            {7'd88,7'd122}:		p = 14'd10736;
            {7'd88,7'd123}:		p = 14'd10824;
            {7'd88,7'd124}:		p = 14'd10912;
            {7'd88,7'd125}:		p = 14'd11000;
            {7'd88,7'd126}:		p = 14'd11088;
            {7'd88,7'd127}:		p = 14'd11176;
            {7'd89,7'd0}:		p = 14'd0;
            {7'd89,7'd1}:		p = 14'd89;
            {7'd89,7'd2}:		p = 14'd178;
            {7'd89,7'd3}:		p = 14'd267;
            {7'd89,7'd4}:		p = 14'd356;
            {7'd89,7'd5}:		p = 14'd445;
            {7'd89,7'd6}:		p = 14'd534;
            {7'd89,7'd7}:		p = 14'd623;
            {7'd89,7'd8}:		p = 14'd712;
            {7'd89,7'd9}:		p = 14'd801;
            {7'd89,7'd10}:		p = 14'd890;
            {7'd89,7'd11}:		p = 14'd979;
            {7'd89,7'd12}:		p = 14'd1068;
            {7'd89,7'd13}:		p = 14'd1157;
            {7'd89,7'd14}:		p = 14'd1246;
            {7'd89,7'd15}:		p = 14'd1335;
            {7'd89,7'd16}:		p = 14'd1424;
            {7'd89,7'd17}:		p = 14'd1513;
            {7'd89,7'd18}:		p = 14'd1602;
            {7'd89,7'd19}:		p = 14'd1691;
            {7'd89,7'd20}:		p = 14'd1780;
            {7'd89,7'd21}:		p = 14'd1869;
            {7'd89,7'd22}:		p = 14'd1958;
            {7'd89,7'd23}:		p = 14'd2047;
            {7'd89,7'd24}:		p = 14'd2136;
            {7'd89,7'd25}:		p = 14'd2225;
            {7'd89,7'd26}:		p = 14'd2314;
            {7'd89,7'd27}:		p = 14'd2403;
            {7'd89,7'd28}:		p = 14'd2492;
            {7'd89,7'd29}:		p = 14'd2581;
            {7'd89,7'd30}:		p = 14'd2670;
            {7'd89,7'd31}:		p = 14'd2759;
            {7'd89,7'd32}:		p = 14'd2848;
            {7'd89,7'd33}:		p = 14'd2937;
            {7'd89,7'd34}:		p = 14'd3026;
            {7'd89,7'd35}:		p = 14'd3115;
            {7'd89,7'd36}:		p = 14'd3204;
            {7'd89,7'd37}:		p = 14'd3293;
            {7'd89,7'd38}:		p = 14'd3382;
            {7'd89,7'd39}:		p = 14'd3471;
            {7'd89,7'd40}:		p = 14'd3560;
            {7'd89,7'd41}:		p = 14'd3649;
            {7'd89,7'd42}:		p = 14'd3738;
            {7'd89,7'd43}:		p = 14'd3827;
            {7'd89,7'd44}:		p = 14'd3916;
            {7'd89,7'd45}:		p = 14'd4005;
            {7'd89,7'd46}:		p = 14'd4094;
            {7'd89,7'd47}:		p = 14'd4183;
            {7'd89,7'd48}:		p = 14'd4272;
            {7'd89,7'd49}:		p = 14'd4361;
            {7'd89,7'd50}:		p = 14'd4450;
            {7'd89,7'd51}:		p = 14'd4539;
            {7'd89,7'd52}:		p = 14'd4628;
            {7'd89,7'd53}:		p = 14'd4717;
            {7'd89,7'd54}:		p = 14'd4806;
            {7'd89,7'd55}:		p = 14'd4895;
            {7'd89,7'd56}:		p = 14'd4984;
            {7'd89,7'd57}:		p = 14'd5073;
            {7'd89,7'd58}:		p = 14'd5162;
            {7'd89,7'd59}:		p = 14'd5251;
            {7'd89,7'd60}:		p = 14'd5340;
            {7'd89,7'd61}:		p = 14'd5429;
            {7'd89,7'd62}:		p = 14'd5518;
            {7'd89,7'd63}:		p = 14'd5607;
            {7'd89,7'd64}:		p = 14'd5696;
            {7'd89,7'd65}:		p = 14'd5785;
            {7'd89,7'd66}:		p = 14'd5874;
            {7'd89,7'd67}:		p = 14'd5963;
            {7'd89,7'd68}:		p = 14'd6052;
            {7'd89,7'd69}:		p = 14'd6141;
            {7'd89,7'd70}:		p = 14'd6230;
            {7'd89,7'd71}:		p = 14'd6319;
            {7'd89,7'd72}:		p = 14'd6408;
            {7'd89,7'd73}:		p = 14'd6497;
            {7'd89,7'd74}:		p = 14'd6586;
            {7'd89,7'd75}:		p = 14'd6675;
            {7'd89,7'd76}:		p = 14'd6764;
            {7'd89,7'd77}:		p = 14'd6853;
            {7'd89,7'd78}:		p = 14'd6942;
            {7'd89,7'd79}:		p = 14'd7031;
            {7'd89,7'd80}:		p = 14'd7120;
            {7'd89,7'd81}:		p = 14'd7209;
            {7'd89,7'd82}:		p = 14'd7298;
            {7'd89,7'd83}:		p = 14'd7387;
            {7'd89,7'd84}:		p = 14'd7476;
            {7'd89,7'd85}:		p = 14'd7565;
            {7'd89,7'd86}:		p = 14'd7654;
            {7'd89,7'd87}:		p = 14'd7743;
            {7'd89,7'd88}:		p = 14'd7832;
            {7'd89,7'd89}:		p = 14'd7921;
            {7'd89,7'd90}:		p = 14'd8010;
            {7'd89,7'd91}:		p = 14'd8099;
            {7'd89,7'd92}:		p = 14'd8188;
            {7'd89,7'd93}:		p = 14'd8277;
            {7'd89,7'd94}:		p = 14'd8366;
            {7'd89,7'd95}:		p = 14'd8455;
            {7'd89,7'd96}:		p = 14'd8544;
            {7'd89,7'd97}:		p = 14'd8633;
            {7'd89,7'd98}:		p = 14'd8722;
            {7'd89,7'd99}:		p = 14'd8811;
            {7'd89,7'd100}:		p = 14'd8900;
            {7'd89,7'd101}:		p = 14'd8989;
            {7'd89,7'd102}:		p = 14'd9078;
            {7'd89,7'd103}:		p = 14'd9167;
            {7'd89,7'd104}:		p = 14'd9256;
            {7'd89,7'd105}:		p = 14'd9345;
            {7'd89,7'd106}:		p = 14'd9434;
            {7'd89,7'd107}:		p = 14'd9523;
            {7'd89,7'd108}:		p = 14'd9612;
            {7'd89,7'd109}:		p = 14'd9701;
            {7'd89,7'd110}:		p = 14'd9790;
            {7'd89,7'd111}:		p = 14'd9879;
            {7'd89,7'd112}:		p = 14'd9968;
            {7'd89,7'd113}:		p = 14'd10057;
            {7'd89,7'd114}:		p = 14'd10146;
            {7'd89,7'd115}:		p = 14'd10235;
            {7'd89,7'd116}:		p = 14'd10324;
            {7'd89,7'd117}:		p = 14'd10413;
            {7'd89,7'd118}:		p = 14'd10502;
            {7'd89,7'd119}:		p = 14'd10591;
            {7'd89,7'd120}:		p = 14'd10680;
            {7'd89,7'd121}:		p = 14'd10769;
            {7'd89,7'd122}:		p = 14'd10858;
            {7'd89,7'd123}:		p = 14'd10947;
            {7'd89,7'd124}:		p = 14'd11036;
            {7'd89,7'd125}:		p = 14'd11125;
            {7'd89,7'd126}:		p = 14'd11214;
            {7'd89,7'd127}:		p = 14'd11303;
            {7'd90,7'd0}:		p = 14'd0;
            {7'd90,7'd1}:		p = 14'd90;
            {7'd90,7'd2}:		p = 14'd180;
            {7'd90,7'd3}:		p = 14'd270;
            {7'd90,7'd4}:		p = 14'd360;
            {7'd90,7'd5}:		p = 14'd450;
            {7'd90,7'd6}:		p = 14'd540;
            {7'd90,7'd7}:		p = 14'd630;
            {7'd90,7'd8}:		p = 14'd720;
            {7'd90,7'd9}:		p = 14'd810;
            {7'd90,7'd10}:		p = 14'd900;
            {7'd90,7'd11}:		p = 14'd990;
            {7'd90,7'd12}:		p = 14'd1080;
            {7'd90,7'd13}:		p = 14'd1170;
            {7'd90,7'd14}:		p = 14'd1260;
            {7'd90,7'd15}:		p = 14'd1350;
            {7'd90,7'd16}:		p = 14'd1440;
            {7'd90,7'd17}:		p = 14'd1530;
            {7'd90,7'd18}:		p = 14'd1620;
            {7'd90,7'd19}:		p = 14'd1710;
            {7'd90,7'd20}:		p = 14'd1800;
            {7'd90,7'd21}:		p = 14'd1890;
            {7'd90,7'd22}:		p = 14'd1980;
            {7'd90,7'd23}:		p = 14'd2070;
            {7'd90,7'd24}:		p = 14'd2160;
            {7'd90,7'd25}:		p = 14'd2250;
            {7'd90,7'd26}:		p = 14'd2340;
            {7'd90,7'd27}:		p = 14'd2430;
            {7'd90,7'd28}:		p = 14'd2520;
            {7'd90,7'd29}:		p = 14'd2610;
            {7'd90,7'd30}:		p = 14'd2700;
            {7'd90,7'd31}:		p = 14'd2790;
            {7'd90,7'd32}:		p = 14'd2880;
            {7'd90,7'd33}:		p = 14'd2970;
            {7'd90,7'd34}:		p = 14'd3060;
            {7'd90,7'd35}:		p = 14'd3150;
            {7'd90,7'd36}:		p = 14'd3240;
            {7'd90,7'd37}:		p = 14'd3330;
            {7'd90,7'd38}:		p = 14'd3420;
            {7'd90,7'd39}:		p = 14'd3510;
            {7'd90,7'd40}:		p = 14'd3600;
            {7'd90,7'd41}:		p = 14'd3690;
            {7'd90,7'd42}:		p = 14'd3780;
            {7'd90,7'd43}:		p = 14'd3870;
            {7'd90,7'd44}:		p = 14'd3960;
            {7'd90,7'd45}:		p = 14'd4050;
            {7'd90,7'd46}:		p = 14'd4140;
            {7'd90,7'd47}:		p = 14'd4230;
            {7'd90,7'd48}:		p = 14'd4320;
            {7'd90,7'd49}:		p = 14'd4410;
            {7'd90,7'd50}:		p = 14'd4500;
            {7'd90,7'd51}:		p = 14'd4590;
            {7'd90,7'd52}:		p = 14'd4680;
            {7'd90,7'd53}:		p = 14'd4770;
            {7'd90,7'd54}:		p = 14'd4860;
            {7'd90,7'd55}:		p = 14'd4950;
            {7'd90,7'd56}:		p = 14'd5040;
            {7'd90,7'd57}:		p = 14'd5130;
            {7'd90,7'd58}:		p = 14'd5220;
            {7'd90,7'd59}:		p = 14'd5310;
            {7'd90,7'd60}:		p = 14'd5400;
            {7'd90,7'd61}:		p = 14'd5490;
            {7'd90,7'd62}:		p = 14'd5580;
            {7'd90,7'd63}:		p = 14'd5670;
            {7'd90,7'd64}:		p = 14'd5760;
            {7'd90,7'd65}:		p = 14'd5850;
            {7'd90,7'd66}:		p = 14'd5940;
            {7'd90,7'd67}:		p = 14'd6030;
            {7'd90,7'd68}:		p = 14'd6120;
            {7'd90,7'd69}:		p = 14'd6210;
            {7'd90,7'd70}:		p = 14'd6300;
            {7'd90,7'd71}:		p = 14'd6390;
            {7'd90,7'd72}:		p = 14'd6480;
            {7'd90,7'd73}:		p = 14'd6570;
            {7'd90,7'd74}:		p = 14'd6660;
            {7'd90,7'd75}:		p = 14'd6750;
            {7'd90,7'd76}:		p = 14'd6840;
            {7'd90,7'd77}:		p = 14'd6930;
            {7'd90,7'd78}:		p = 14'd7020;
            {7'd90,7'd79}:		p = 14'd7110;
            {7'd90,7'd80}:		p = 14'd7200;
            {7'd90,7'd81}:		p = 14'd7290;
            {7'd90,7'd82}:		p = 14'd7380;
            {7'd90,7'd83}:		p = 14'd7470;
            {7'd90,7'd84}:		p = 14'd7560;
            {7'd90,7'd85}:		p = 14'd7650;
            {7'd90,7'd86}:		p = 14'd7740;
            {7'd90,7'd87}:		p = 14'd7830;
            {7'd90,7'd88}:		p = 14'd7920;
            {7'd90,7'd89}:		p = 14'd8010;
            {7'd90,7'd90}:		p = 14'd8100;
            {7'd90,7'd91}:		p = 14'd8190;
            {7'd90,7'd92}:		p = 14'd8280;
            {7'd90,7'd93}:		p = 14'd8370;
            {7'd90,7'd94}:		p = 14'd8460;
            {7'd90,7'd95}:		p = 14'd8550;
            {7'd90,7'd96}:		p = 14'd8640;
            {7'd90,7'd97}:		p = 14'd8730;
            {7'd90,7'd98}:		p = 14'd8820;
            {7'd90,7'd99}:		p = 14'd8910;
            {7'd90,7'd100}:		p = 14'd9000;
            {7'd90,7'd101}:		p = 14'd9090;
            {7'd90,7'd102}:		p = 14'd9180;
            {7'd90,7'd103}:		p = 14'd9270;
            {7'd90,7'd104}:		p = 14'd9360;
            {7'd90,7'd105}:		p = 14'd9450;
            {7'd90,7'd106}:		p = 14'd9540;
            {7'd90,7'd107}:		p = 14'd9630;
            {7'd90,7'd108}:		p = 14'd9720;
            {7'd90,7'd109}:		p = 14'd9810;
            {7'd90,7'd110}:		p = 14'd9900;
            {7'd90,7'd111}:		p = 14'd9990;
            {7'd90,7'd112}:		p = 14'd10080;
            {7'd90,7'd113}:		p = 14'd10170;
            {7'd90,7'd114}:		p = 14'd10260;
            {7'd90,7'd115}:		p = 14'd10350;
            {7'd90,7'd116}:		p = 14'd10440;
            {7'd90,7'd117}:		p = 14'd10530;
            {7'd90,7'd118}:		p = 14'd10620;
            {7'd90,7'd119}:		p = 14'd10710;
            {7'd90,7'd120}:		p = 14'd10800;
            {7'd90,7'd121}:		p = 14'd10890;
            {7'd90,7'd122}:		p = 14'd10980;
            {7'd90,7'd123}:		p = 14'd11070;
            {7'd90,7'd124}:		p = 14'd11160;
            {7'd90,7'd125}:		p = 14'd11250;
            {7'd90,7'd126}:		p = 14'd11340;
            {7'd90,7'd127}:		p = 14'd11430;
            {7'd91,7'd0}:		p = 14'd0;
            {7'd91,7'd1}:		p = 14'd91;
            {7'd91,7'd2}:		p = 14'd182;
            {7'd91,7'd3}:		p = 14'd273;
            {7'd91,7'd4}:		p = 14'd364;
            {7'd91,7'd5}:		p = 14'd455;
            {7'd91,7'd6}:		p = 14'd546;
            {7'd91,7'd7}:		p = 14'd637;
            {7'd91,7'd8}:		p = 14'd728;
            {7'd91,7'd9}:		p = 14'd819;
            {7'd91,7'd10}:		p = 14'd910;
            {7'd91,7'd11}:		p = 14'd1001;
            {7'd91,7'd12}:		p = 14'd1092;
            {7'd91,7'd13}:		p = 14'd1183;
            {7'd91,7'd14}:		p = 14'd1274;
            {7'd91,7'd15}:		p = 14'd1365;
            {7'd91,7'd16}:		p = 14'd1456;
            {7'd91,7'd17}:		p = 14'd1547;
            {7'd91,7'd18}:		p = 14'd1638;
            {7'd91,7'd19}:		p = 14'd1729;
            {7'd91,7'd20}:		p = 14'd1820;
            {7'd91,7'd21}:		p = 14'd1911;
            {7'd91,7'd22}:		p = 14'd2002;
            {7'd91,7'd23}:		p = 14'd2093;
            {7'd91,7'd24}:		p = 14'd2184;
            {7'd91,7'd25}:		p = 14'd2275;
            {7'd91,7'd26}:		p = 14'd2366;
            {7'd91,7'd27}:		p = 14'd2457;
            {7'd91,7'd28}:		p = 14'd2548;
            {7'd91,7'd29}:		p = 14'd2639;
            {7'd91,7'd30}:		p = 14'd2730;
            {7'd91,7'd31}:		p = 14'd2821;
            {7'd91,7'd32}:		p = 14'd2912;
            {7'd91,7'd33}:		p = 14'd3003;
            {7'd91,7'd34}:		p = 14'd3094;
            {7'd91,7'd35}:		p = 14'd3185;
            {7'd91,7'd36}:		p = 14'd3276;
            {7'd91,7'd37}:		p = 14'd3367;
            {7'd91,7'd38}:		p = 14'd3458;
            {7'd91,7'd39}:		p = 14'd3549;
            {7'd91,7'd40}:		p = 14'd3640;
            {7'd91,7'd41}:		p = 14'd3731;
            {7'd91,7'd42}:		p = 14'd3822;
            {7'd91,7'd43}:		p = 14'd3913;
            {7'd91,7'd44}:		p = 14'd4004;
            {7'd91,7'd45}:		p = 14'd4095;
            {7'd91,7'd46}:		p = 14'd4186;
            {7'd91,7'd47}:		p = 14'd4277;
            {7'd91,7'd48}:		p = 14'd4368;
            {7'd91,7'd49}:		p = 14'd4459;
            {7'd91,7'd50}:		p = 14'd4550;
            {7'd91,7'd51}:		p = 14'd4641;
            {7'd91,7'd52}:		p = 14'd4732;
            {7'd91,7'd53}:		p = 14'd4823;
            {7'd91,7'd54}:		p = 14'd4914;
            {7'd91,7'd55}:		p = 14'd5005;
            {7'd91,7'd56}:		p = 14'd5096;
            {7'd91,7'd57}:		p = 14'd5187;
            {7'd91,7'd58}:		p = 14'd5278;
            {7'd91,7'd59}:		p = 14'd5369;
            {7'd91,7'd60}:		p = 14'd5460;
            {7'd91,7'd61}:		p = 14'd5551;
            {7'd91,7'd62}:		p = 14'd5642;
            {7'd91,7'd63}:		p = 14'd5733;
            {7'd91,7'd64}:		p = 14'd5824;
            {7'd91,7'd65}:		p = 14'd5915;
            {7'd91,7'd66}:		p = 14'd6006;
            {7'd91,7'd67}:		p = 14'd6097;
            {7'd91,7'd68}:		p = 14'd6188;
            {7'd91,7'd69}:		p = 14'd6279;
            {7'd91,7'd70}:		p = 14'd6370;
            {7'd91,7'd71}:		p = 14'd6461;
            {7'd91,7'd72}:		p = 14'd6552;
            {7'd91,7'd73}:		p = 14'd6643;
            {7'd91,7'd74}:		p = 14'd6734;
            {7'd91,7'd75}:		p = 14'd6825;
            {7'd91,7'd76}:		p = 14'd6916;
            {7'd91,7'd77}:		p = 14'd7007;
            {7'd91,7'd78}:		p = 14'd7098;
            {7'd91,7'd79}:		p = 14'd7189;
            {7'd91,7'd80}:		p = 14'd7280;
            {7'd91,7'd81}:		p = 14'd7371;
            {7'd91,7'd82}:		p = 14'd7462;
            {7'd91,7'd83}:		p = 14'd7553;
            {7'd91,7'd84}:		p = 14'd7644;
            {7'd91,7'd85}:		p = 14'd7735;
            {7'd91,7'd86}:		p = 14'd7826;
            {7'd91,7'd87}:		p = 14'd7917;
            {7'd91,7'd88}:		p = 14'd8008;
            {7'd91,7'd89}:		p = 14'd8099;
            {7'd91,7'd90}:		p = 14'd8190;
            {7'd91,7'd91}:		p = 14'd8281;
            {7'd91,7'd92}:		p = 14'd8372;
            {7'd91,7'd93}:		p = 14'd8463;
            {7'd91,7'd94}:		p = 14'd8554;
            {7'd91,7'd95}:		p = 14'd8645;
            {7'd91,7'd96}:		p = 14'd8736;
            {7'd91,7'd97}:		p = 14'd8827;
            {7'd91,7'd98}:		p = 14'd8918;
            {7'd91,7'd99}:		p = 14'd9009;
            {7'd91,7'd100}:		p = 14'd9100;
            {7'd91,7'd101}:		p = 14'd9191;
            {7'd91,7'd102}:		p = 14'd9282;
            {7'd91,7'd103}:		p = 14'd9373;
            {7'd91,7'd104}:		p = 14'd9464;
            {7'd91,7'd105}:		p = 14'd9555;
            {7'd91,7'd106}:		p = 14'd9646;
            {7'd91,7'd107}:		p = 14'd9737;
            {7'd91,7'd108}:		p = 14'd9828;
            {7'd91,7'd109}:		p = 14'd9919;
            {7'd91,7'd110}:		p = 14'd10010;
            {7'd91,7'd111}:		p = 14'd10101;
            {7'd91,7'd112}:		p = 14'd10192;
            {7'd91,7'd113}:		p = 14'd10283;
            {7'd91,7'd114}:		p = 14'd10374;
            {7'd91,7'd115}:		p = 14'd10465;
            {7'd91,7'd116}:		p = 14'd10556;
            {7'd91,7'd117}:		p = 14'd10647;
            {7'd91,7'd118}:		p = 14'd10738;
            {7'd91,7'd119}:		p = 14'd10829;
            {7'd91,7'd120}:		p = 14'd10920;
            {7'd91,7'd121}:		p = 14'd11011;
            {7'd91,7'd122}:		p = 14'd11102;
            {7'd91,7'd123}:		p = 14'd11193;
            {7'd91,7'd124}:		p = 14'd11284;
            {7'd91,7'd125}:		p = 14'd11375;
            {7'd91,7'd126}:		p = 14'd11466;
            {7'd91,7'd127}:		p = 14'd11557;
            {7'd92,7'd0}:		p = 14'd0;
            {7'd92,7'd1}:		p = 14'd92;
            {7'd92,7'd2}:		p = 14'd184;
            {7'd92,7'd3}:		p = 14'd276;
            {7'd92,7'd4}:		p = 14'd368;
            {7'd92,7'd5}:		p = 14'd460;
            {7'd92,7'd6}:		p = 14'd552;
            {7'd92,7'd7}:		p = 14'd644;
            {7'd92,7'd8}:		p = 14'd736;
            {7'd92,7'd9}:		p = 14'd828;
            {7'd92,7'd10}:		p = 14'd920;
            {7'd92,7'd11}:		p = 14'd1012;
            {7'd92,7'd12}:		p = 14'd1104;
            {7'd92,7'd13}:		p = 14'd1196;
            {7'd92,7'd14}:		p = 14'd1288;
            {7'd92,7'd15}:		p = 14'd1380;
            {7'd92,7'd16}:		p = 14'd1472;
            {7'd92,7'd17}:		p = 14'd1564;
            {7'd92,7'd18}:		p = 14'd1656;
            {7'd92,7'd19}:		p = 14'd1748;
            {7'd92,7'd20}:		p = 14'd1840;
            {7'd92,7'd21}:		p = 14'd1932;
            {7'd92,7'd22}:		p = 14'd2024;
            {7'd92,7'd23}:		p = 14'd2116;
            {7'd92,7'd24}:		p = 14'd2208;
            {7'd92,7'd25}:		p = 14'd2300;
            {7'd92,7'd26}:		p = 14'd2392;
            {7'd92,7'd27}:		p = 14'd2484;
            {7'd92,7'd28}:		p = 14'd2576;
            {7'd92,7'd29}:		p = 14'd2668;
            {7'd92,7'd30}:		p = 14'd2760;
            {7'd92,7'd31}:		p = 14'd2852;
            {7'd92,7'd32}:		p = 14'd2944;
            {7'd92,7'd33}:		p = 14'd3036;
            {7'd92,7'd34}:		p = 14'd3128;
            {7'd92,7'd35}:		p = 14'd3220;
            {7'd92,7'd36}:		p = 14'd3312;
            {7'd92,7'd37}:		p = 14'd3404;
            {7'd92,7'd38}:		p = 14'd3496;
            {7'd92,7'd39}:		p = 14'd3588;
            {7'd92,7'd40}:		p = 14'd3680;
            {7'd92,7'd41}:		p = 14'd3772;
            {7'd92,7'd42}:		p = 14'd3864;
            {7'd92,7'd43}:		p = 14'd3956;
            {7'd92,7'd44}:		p = 14'd4048;
            {7'd92,7'd45}:		p = 14'd4140;
            {7'd92,7'd46}:		p = 14'd4232;
            {7'd92,7'd47}:		p = 14'd4324;
            {7'd92,7'd48}:		p = 14'd4416;
            {7'd92,7'd49}:		p = 14'd4508;
            {7'd92,7'd50}:		p = 14'd4600;
            {7'd92,7'd51}:		p = 14'd4692;
            {7'd92,7'd52}:		p = 14'd4784;
            {7'd92,7'd53}:		p = 14'd4876;
            {7'd92,7'd54}:		p = 14'd4968;
            {7'd92,7'd55}:		p = 14'd5060;
            {7'd92,7'd56}:		p = 14'd5152;
            {7'd92,7'd57}:		p = 14'd5244;
            {7'd92,7'd58}:		p = 14'd5336;
            {7'd92,7'd59}:		p = 14'd5428;
            {7'd92,7'd60}:		p = 14'd5520;
            {7'd92,7'd61}:		p = 14'd5612;
            {7'd92,7'd62}:		p = 14'd5704;
            {7'd92,7'd63}:		p = 14'd5796;
            {7'd92,7'd64}:		p = 14'd5888;
            {7'd92,7'd65}:		p = 14'd5980;
            {7'd92,7'd66}:		p = 14'd6072;
            {7'd92,7'd67}:		p = 14'd6164;
            {7'd92,7'd68}:		p = 14'd6256;
            {7'd92,7'd69}:		p = 14'd6348;
            {7'd92,7'd70}:		p = 14'd6440;
            {7'd92,7'd71}:		p = 14'd6532;
            {7'd92,7'd72}:		p = 14'd6624;
            {7'd92,7'd73}:		p = 14'd6716;
            {7'd92,7'd74}:		p = 14'd6808;
            {7'd92,7'd75}:		p = 14'd6900;
            {7'd92,7'd76}:		p = 14'd6992;
            {7'd92,7'd77}:		p = 14'd7084;
            {7'd92,7'd78}:		p = 14'd7176;
            {7'd92,7'd79}:		p = 14'd7268;
            {7'd92,7'd80}:		p = 14'd7360;
            {7'd92,7'd81}:		p = 14'd7452;
            {7'd92,7'd82}:		p = 14'd7544;
            {7'd92,7'd83}:		p = 14'd7636;
            {7'd92,7'd84}:		p = 14'd7728;
            {7'd92,7'd85}:		p = 14'd7820;
            {7'd92,7'd86}:		p = 14'd7912;
            {7'd92,7'd87}:		p = 14'd8004;
            {7'd92,7'd88}:		p = 14'd8096;
            {7'd92,7'd89}:		p = 14'd8188;
            {7'd92,7'd90}:		p = 14'd8280;
            {7'd92,7'd91}:		p = 14'd8372;
            {7'd92,7'd92}:		p = 14'd8464;
            {7'd92,7'd93}:		p = 14'd8556;
            {7'd92,7'd94}:		p = 14'd8648;
            {7'd92,7'd95}:		p = 14'd8740;
            {7'd92,7'd96}:		p = 14'd8832;
            {7'd92,7'd97}:		p = 14'd8924;
            {7'd92,7'd98}:		p = 14'd9016;
            {7'd92,7'd99}:		p = 14'd9108;
            {7'd92,7'd100}:		p = 14'd9200;
            {7'd92,7'd101}:		p = 14'd9292;
            {7'd92,7'd102}:		p = 14'd9384;
            {7'd92,7'd103}:		p = 14'd9476;
            {7'd92,7'd104}:		p = 14'd9568;
            {7'd92,7'd105}:		p = 14'd9660;
            {7'd92,7'd106}:		p = 14'd9752;
            {7'd92,7'd107}:		p = 14'd9844;
            {7'd92,7'd108}:		p = 14'd9936;
            {7'd92,7'd109}:		p = 14'd10028;
            {7'd92,7'd110}:		p = 14'd10120;
            {7'd92,7'd111}:		p = 14'd10212;
            {7'd92,7'd112}:		p = 14'd10304;
            {7'd92,7'd113}:		p = 14'd10396;
            {7'd92,7'd114}:		p = 14'd10488;
            {7'd92,7'd115}:		p = 14'd10580;
            {7'd92,7'd116}:		p = 14'd10672;
            {7'd92,7'd117}:		p = 14'd10764;
            {7'd92,7'd118}:		p = 14'd10856;
            {7'd92,7'd119}:		p = 14'd10948;
            {7'd92,7'd120}:		p = 14'd11040;
            {7'd92,7'd121}:		p = 14'd11132;
            {7'd92,7'd122}:		p = 14'd11224;
            {7'd92,7'd123}:		p = 14'd11316;
            {7'd92,7'd124}:		p = 14'd11408;
            {7'd92,7'd125}:		p = 14'd11500;
            {7'd92,7'd126}:		p = 14'd11592;
            {7'd92,7'd127}:		p = 14'd11684;
            {7'd93,7'd0}:		p = 14'd0;
            {7'd93,7'd1}:		p = 14'd93;
            {7'd93,7'd2}:		p = 14'd186;
            {7'd93,7'd3}:		p = 14'd279;
            {7'd93,7'd4}:		p = 14'd372;
            {7'd93,7'd5}:		p = 14'd465;
            {7'd93,7'd6}:		p = 14'd558;
            {7'd93,7'd7}:		p = 14'd651;
            {7'd93,7'd8}:		p = 14'd744;
            {7'd93,7'd9}:		p = 14'd837;
            {7'd93,7'd10}:		p = 14'd930;
            {7'd93,7'd11}:		p = 14'd1023;
            {7'd93,7'd12}:		p = 14'd1116;
            {7'd93,7'd13}:		p = 14'd1209;
            {7'd93,7'd14}:		p = 14'd1302;
            {7'd93,7'd15}:		p = 14'd1395;
            {7'd93,7'd16}:		p = 14'd1488;
            {7'd93,7'd17}:		p = 14'd1581;
            {7'd93,7'd18}:		p = 14'd1674;
            {7'd93,7'd19}:		p = 14'd1767;
            {7'd93,7'd20}:		p = 14'd1860;
            {7'd93,7'd21}:		p = 14'd1953;
            {7'd93,7'd22}:		p = 14'd2046;
            {7'd93,7'd23}:		p = 14'd2139;
            {7'd93,7'd24}:		p = 14'd2232;
            {7'd93,7'd25}:		p = 14'd2325;
            {7'd93,7'd26}:		p = 14'd2418;
            {7'd93,7'd27}:		p = 14'd2511;
            {7'd93,7'd28}:		p = 14'd2604;
            {7'd93,7'd29}:		p = 14'd2697;
            {7'd93,7'd30}:		p = 14'd2790;
            {7'd93,7'd31}:		p = 14'd2883;
            {7'd93,7'd32}:		p = 14'd2976;
            {7'd93,7'd33}:		p = 14'd3069;
            {7'd93,7'd34}:		p = 14'd3162;
            {7'd93,7'd35}:		p = 14'd3255;
            {7'd93,7'd36}:		p = 14'd3348;
            {7'd93,7'd37}:		p = 14'd3441;
            {7'd93,7'd38}:		p = 14'd3534;
            {7'd93,7'd39}:		p = 14'd3627;
            {7'd93,7'd40}:		p = 14'd3720;
            {7'd93,7'd41}:		p = 14'd3813;
            {7'd93,7'd42}:		p = 14'd3906;
            {7'd93,7'd43}:		p = 14'd3999;
            {7'd93,7'd44}:		p = 14'd4092;
            {7'd93,7'd45}:		p = 14'd4185;
            {7'd93,7'd46}:		p = 14'd4278;
            {7'd93,7'd47}:		p = 14'd4371;
            {7'd93,7'd48}:		p = 14'd4464;
            {7'd93,7'd49}:		p = 14'd4557;
            {7'd93,7'd50}:		p = 14'd4650;
            {7'd93,7'd51}:		p = 14'd4743;
            {7'd93,7'd52}:		p = 14'd4836;
            {7'd93,7'd53}:		p = 14'd4929;
            {7'd93,7'd54}:		p = 14'd5022;
            {7'd93,7'd55}:		p = 14'd5115;
            {7'd93,7'd56}:		p = 14'd5208;
            {7'd93,7'd57}:		p = 14'd5301;
            {7'd93,7'd58}:		p = 14'd5394;
            {7'd93,7'd59}:		p = 14'd5487;
            {7'd93,7'd60}:		p = 14'd5580;
            {7'd93,7'd61}:		p = 14'd5673;
            {7'd93,7'd62}:		p = 14'd5766;
            {7'd93,7'd63}:		p = 14'd5859;
            {7'd93,7'd64}:		p = 14'd5952;
            {7'd93,7'd65}:		p = 14'd6045;
            {7'd93,7'd66}:		p = 14'd6138;
            {7'd93,7'd67}:		p = 14'd6231;
            {7'd93,7'd68}:		p = 14'd6324;
            {7'd93,7'd69}:		p = 14'd6417;
            {7'd93,7'd70}:		p = 14'd6510;
            {7'd93,7'd71}:		p = 14'd6603;
            {7'd93,7'd72}:		p = 14'd6696;
            {7'd93,7'd73}:		p = 14'd6789;
            {7'd93,7'd74}:		p = 14'd6882;
            {7'd93,7'd75}:		p = 14'd6975;
            {7'd93,7'd76}:		p = 14'd7068;
            {7'd93,7'd77}:		p = 14'd7161;
            {7'd93,7'd78}:		p = 14'd7254;
            {7'd93,7'd79}:		p = 14'd7347;
            {7'd93,7'd80}:		p = 14'd7440;
            {7'd93,7'd81}:		p = 14'd7533;
            {7'd93,7'd82}:		p = 14'd7626;
            {7'd93,7'd83}:		p = 14'd7719;
            {7'd93,7'd84}:		p = 14'd7812;
            {7'd93,7'd85}:		p = 14'd7905;
            {7'd93,7'd86}:		p = 14'd7998;
            {7'd93,7'd87}:		p = 14'd8091;
            {7'd93,7'd88}:		p = 14'd8184;
            {7'd93,7'd89}:		p = 14'd8277;
            {7'd93,7'd90}:		p = 14'd8370;
            {7'd93,7'd91}:		p = 14'd8463;
            {7'd93,7'd92}:		p = 14'd8556;
            {7'd93,7'd93}:		p = 14'd8649;
            {7'd93,7'd94}:		p = 14'd8742;
            {7'd93,7'd95}:		p = 14'd8835;
            {7'd93,7'd96}:		p = 14'd8928;
            {7'd93,7'd97}:		p = 14'd9021;
            {7'd93,7'd98}:		p = 14'd9114;
            {7'd93,7'd99}:		p = 14'd9207;
            {7'd93,7'd100}:		p = 14'd9300;
            {7'd93,7'd101}:		p = 14'd9393;
            {7'd93,7'd102}:		p = 14'd9486;
            {7'd93,7'd103}:		p = 14'd9579;
            {7'd93,7'd104}:		p = 14'd9672;
            {7'd93,7'd105}:		p = 14'd9765;
            {7'd93,7'd106}:		p = 14'd9858;
            {7'd93,7'd107}:		p = 14'd9951;
            {7'd93,7'd108}:		p = 14'd10044;
            {7'd93,7'd109}:		p = 14'd10137;
            {7'd93,7'd110}:		p = 14'd10230;
            {7'd93,7'd111}:		p = 14'd10323;
            {7'd93,7'd112}:		p = 14'd10416;
            {7'd93,7'd113}:		p = 14'd10509;
            {7'd93,7'd114}:		p = 14'd10602;
            {7'd93,7'd115}:		p = 14'd10695;
            {7'd93,7'd116}:		p = 14'd10788;
            {7'd93,7'd117}:		p = 14'd10881;
            {7'd93,7'd118}:		p = 14'd10974;
            {7'd93,7'd119}:		p = 14'd11067;
            {7'd93,7'd120}:		p = 14'd11160;
            {7'd93,7'd121}:		p = 14'd11253;
            {7'd93,7'd122}:		p = 14'd11346;
            {7'd93,7'd123}:		p = 14'd11439;
            {7'd93,7'd124}:		p = 14'd11532;
            {7'd93,7'd125}:		p = 14'd11625;
            {7'd93,7'd126}:		p = 14'd11718;
            {7'd93,7'd127}:		p = 14'd11811;
            {7'd94,7'd0}:		p = 14'd0;
            {7'd94,7'd1}:		p = 14'd94;
            {7'd94,7'd2}:		p = 14'd188;
            {7'd94,7'd3}:		p = 14'd282;
            {7'd94,7'd4}:		p = 14'd376;
            {7'd94,7'd5}:		p = 14'd470;
            {7'd94,7'd6}:		p = 14'd564;
            {7'd94,7'd7}:		p = 14'd658;
            {7'd94,7'd8}:		p = 14'd752;
            {7'd94,7'd9}:		p = 14'd846;
            {7'd94,7'd10}:		p = 14'd940;
            {7'd94,7'd11}:		p = 14'd1034;
            {7'd94,7'd12}:		p = 14'd1128;
            {7'd94,7'd13}:		p = 14'd1222;
            {7'd94,7'd14}:		p = 14'd1316;
            {7'd94,7'd15}:		p = 14'd1410;
            {7'd94,7'd16}:		p = 14'd1504;
            {7'd94,7'd17}:		p = 14'd1598;
            {7'd94,7'd18}:		p = 14'd1692;
            {7'd94,7'd19}:		p = 14'd1786;
            {7'd94,7'd20}:		p = 14'd1880;
            {7'd94,7'd21}:		p = 14'd1974;
            {7'd94,7'd22}:		p = 14'd2068;
            {7'd94,7'd23}:		p = 14'd2162;
            {7'd94,7'd24}:		p = 14'd2256;
            {7'd94,7'd25}:		p = 14'd2350;
            {7'd94,7'd26}:		p = 14'd2444;
            {7'd94,7'd27}:		p = 14'd2538;
            {7'd94,7'd28}:		p = 14'd2632;
            {7'd94,7'd29}:		p = 14'd2726;
            {7'd94,7'd30}:		p = 14'd2820;
            {7'd94,7'd31}:		p = 14'd2914;
            {7'd94,7'd32}:		p = 14'd3008;
            {7'd94,7'd33}:		p = 14'd3102;
            {7'd94,7'd34}:		p = 14'd3196;
            {7'd94,7'd35}:		p = 14'd3290;
            {7'd94,7'd36}:		p = 14'd3384;
            {7'd94,7'd37}:		p = 14'd3478;
            {7'd94,7'd38}:		p = 14'd3572;
            {7'd94,7'd39}:		p = 14'd3666;
            {7'd94,7'd40}:		p = 14'd3760;
            {7'd94,7'd41}:		p = 14'd3854;
            {7'd94,7'd42}:		p = 14'd3948;
            {7'd94,7'd43}:		p = 14'd4042;
            {7'd94,7'd44}:		p = 14'd4136;
            {7'd94,7'd45}:		p = 14'd4230;
            {7'd94,7'd46}:		p = 14'd4324;
            {7'd94,7'd47}:		p = 14'd4418;
            {7'd94,7'd48}:		p = 14'd4512;
            {7'd94,7'd49}:		p = 14'd4606;
            {7'd94,7'd50}:		p = 14'd4700;
            {7'd94,7'd51}:		p = 14'd4794;
            {7'd94,7'd52}:		p = 14'd4888;
            {7'd94,7'd53}:		p = 14'd4982;
            {7'd94,7'd54}:		p = 14'd5076;
            {7'd94,7'd55}:		p = 14'd5170;
            {7'd94,7'd56}:		p = 14'd5264;
            {7'd94,7'd57}:		p = 14'd5358;
            {7'd94,7'd58}:		p = 14'd5452;
            {7'd94,7'd59}:		p = 14'd5546;
            {7'd94,7'd60}:		p = 14'd5640;
            {7'd94,7'd61}:		p = 14'd5734;
            {7'd94,7'd62}:		p = 14'd5828;
            {7'd94,7'd63}:		p = 14'd5922;
            {7'd94,7'd64}:		p = 14'd6016;
            {7'd94,7'd65}:		p = 14'd6110;
            {7'd94,7'd66}:		p = 14'd6204;
            {7'd94,7'd67}:		p = 14'd6298;
            {7'd94,7'd68}:		p = 14'd6392;
            {7'd94,7'd69}:		p = 14'd6486;
            {7'd94,7'd70}:		p = 14'd6580;
            {7'd94,7'd71}:		p = 14'd6674;
            {7'd94,7'd72}:		p = 14'd6768;
            {7'd94,7'd73}:		p = 14'd6862;
            {7'd94,7'd74}:		p = 14'd6956;
            {7'd94,7'd75}:		p = 14'd7050;
            {7'd94,7'd76}:		p = 14'd7144;
            {7'd94,7'd77}:		p = 14'd7238;
            {7'd94,7'd78}:		p = 14'd7332;
            {7'd94,7'd79}:		p = 14'd7426;
            {7'd94,7'd80}:		p = 14'd7520;
            {7'd94,7'd81}:		p = 14'd7614;
            {7'd94,7'd82}:		p = 14'd7708;
            {7'd94,7'd83}:		p = 14'd7802;
            {7'd94,7'd84}:		p = 14'd7896;
            {7'd94,7'd85}:		p = 14'd7990;
            {7'd94,7'd86}:		p = 14'd8084;
            {7'd94,7'd87}:		p = 14'd8178;
            {7'd94,7'd88}:		p = 14'd8272;
            {7'd94,7'd89}:		p = 14'd8366;
            {7'd94,7'd90}:		p = 14'd8460;
            {7'd94,7'd91}:		p = 14'd8554;
            {7'd94,7'd92}:		p = 14'd8648;
            {7'd94,7'd93}:		p = 14'd8742;
            {7'd94,7'd94}:		p = 14'd8836;
            {7'd94,7'd95}:		p = 14'd8930;
            {7'd94,7'd96}:		p = 14'd9024;
            {7'd94,7'd97}:		p = 14'd9118;
            {7'd94,7'd98}:		p = 14'd9212;
            {7'd94,7'd99}:		p = 14'd9306;
            {7'd94,7'd100}:		p = 14'd9400;
            {7'd94,7'd101}:		p = 14'd9494;
            {7'd94,7'd102}:		p = 14'd9588;
            {7'd94,7'd103}:		p = 14'd9682;
            {7'd94,7'd104}:		p = 14'd9776;
            {7'd94,7'd105}:		p = 14'd9870;
            {7'd94,7'd106}:		p = 14'd9964;
            {7'd94,7'd107}:		p = 14'd10058;
            {7'd94,7'd108}:		p = 14'd10152;
            {7'd94,7'd109}:		p = 14'd10246;
            {7'd94,7'd110}:		p = 14'd10340;
            {7'd94,7'd111}:		p = 14'd10434;
            {7'd94,7'd112}:		p = 14'd10528;
            {7'd94,7'd113}:		p = 14'd10622;
            {7'd94,7'd114}:		p = 14'd10716;
            {7'd94,7'd115}:		p = 14'd10810;
            {7'd94,7'd116}:		p = 14'd10904;
            {7'd94,7'd117}:		p = 14'd10998;
            {7'd94,7'd118}:		p = 14'd11092;
            {7'd94,7'd119}:		p = 14'd11186;
            {7'd94,7'd120}:		p = 14'd11280;
            {7'd94,7'd121}:		p = 14'd11374;
            {7'd94,7'd122}:		p = 14'd11468;
            {7'd94,7'd123}:		p = 14'd11562;
            {7'd94,7'd124}:		p = 14'd11656;
            {7'd94,7'd125}:		p = 14'd11750;
            {7'd94,7'd126}:		p = 14'd11844;
            {7'd94,7'd127}:		p = 14'd11938;
            {7'd95,7'd0}:		p = 14'd0;
            {7'd95,7'd1}:		p = 14'd95;
            {7'd95,7'd2}:		p = 14'd190;
            {7'd95,7'd3}:		p = 14'd285;
            {7'd95,7'd4}:		p = 14'd380;
            {7'd95,7'd5}:		p = 14'd475;
            {7'd95,7'd6}:		p = 14'd570;
            {7'd95,7'd7}:		p = 14'd665;
            {7'd95,7'd8}:		p = 14'd760;
            {7'd95,7'd9}:		p = 14'd855;
            {7'd95,7'd10}:		p = 14'd950;
            {7'd95,7'd11}:		p = 14'd1045;
            {7'd95,7'd12}:		p = 14'd1140;
            {7'd95,7'd13}:		p = 14'd1235;
            {7'd95,7'd14}:		p = 14'd1330;
            {7'd95,7'd15}:		p = 14'd1425;
            {7'd95,7'd16}:		p = 14'd1520;
            {7'd95,7'd17}:		p = 14'd1615;
            {7'd95,7'd18}:		p = 14'd1710;
            {7'd95,7'd19}:		p = 14'd1805;
            {7'd95,7'd20}:		p = 14'd1900;
            {7'd95,7'd21}:		p = 14'd1995;
            {7'd95,7'd22}:		p = 14'd2090;
            {7'd95,7'd23}:		p = 14'd2185;
            {7'd95,7'd24}:		p = 14'd2280;
            {7'd95,7'd25}:		p = 14'd2375;
            {7'd95,7'd26}:		p = 14'd2470;
            {7'd95,7'd27}:		p = 14'd2565;
            {7'd95,7'd28}:		p = 14'd2660;
            {7'd95,7'd29}:		p = 14'd2755;
            {7'd95,7'd30}:		p = 14'd2850;
            {7'd95,7'd31}:		p = 14'd2945;
            {7'd95,7'd32}:		p = 14'd3040;
            {7'd95,7'd33}:		p = 14'd3135;
            {7'd95,7'd34}:		p = 14'd3230;
            {7'd95,7'd35}:		p = 14'd3325;
            {7'd95,7'd36}:		p = 14'd3420;
            {7'd95,7'd37}:		p = 14'd3515;
            {7'd95,7'd38}:		p = 14'd3610;
            {7'd95,7'd39}:		p = 14'd3705;
            {7'd95,7'd40}:		p = 14'd3800;
            {7'd95,7'd41}:		p = 14'd3895;
            {7'd95,7'd42}:		p = 14'd3990;
            {7'd95,7'd43}:		p = 14'd4085;
            {7'd95,7'd44}:		p = 14'd4180;
            {7'd95,7'd45}:		p = 14'd4275;
            {7'd95,7'd46}:		p = 14'd4370;
            {7'd95,7'd47}:		p = 14'd4465;
            {7'd95,7'd48}:		p = 14'd4560;
            {7'd95,7'd49}:		p = 14'd4655;
            {7'd95,7'd50}:		p = 14'd4750;
            {7'd95,7'd51}:		p = 14'd4845;
            {7'd95,7'd52}:		p = 14'd4940;
            {7'd95,7'd53}:		p = 14'd5035;
            {7'd95,7'd54}:		p = 14'd5130;
            {7'd95,7'd55}:		p = 14'd5225;
            {7'd95,7'd56}:		p = 14'd5320;
            {7'd95,7'd57}:		p = 14'd5415;
            {7'd95,7'd58}:		p = 14'd5510;
            {7'd95,7'd59}:		p = 14'd5605;
            {7'd95,7'd60}:		p = 14'd5700;
            {7'd95,7'd61}:		p = 14'd5795;
            {7'd95,7'd62}:		p = 14'd5890;
            {7'd95,7'd63}:		p = 14'd5985;
            {7'd95,7'd64}:		p = 14'd6080;
            {7'd95,7'd65}:		p = 14'd6175;
            {7'd95,7'd66}:		p = 14'd6270;
            {7'd95,7'd67}:		p = 14'd6365;
            {7'd95,7'd68}:		p = 14'd6460;
            {7'd95,7'd69}:		p = 14'd6555;
            {7'd95,7'd70}:		p = 14'd6650;
            {7'd95,7'd71}:		p = 14'd6745;
            {7'd95,7'd72}:		p = 14'd6840;
            {7'd95,7'd73}:		p = 14'd6935;
            {7'd95,7'd74}:		p = 14'd7030;
            {7'd95,7'd75}:		p = 14'd7125;
            {7'd95,7'd76}:		p = 14'd7220;
            {7'd95,7'd77}:		p = 14'd7315;
            {7'd95,7'd78}:		p = 14'd7410;
            {7'd95,7'd79}:		p = 14'd7505;
            {7'd95,7'd80}:		p = 14'd7600;
            {7'd95,7'd81}:		p = 14'd7695;
            {7'd95,7'd82}:		p = 14'd7790;
            {7'd95,7'd83}:		p = 14'd7885;
            {7'd95,7'd84}:		p = 14'd7980;
            {7'd95,7'd85}:		p = 14'd8075;
            {7'd95,7'd86}:		p = 14'd8170;
            {7'd95,7'd87}:		p = 14'd8265;
            {7'd95,7'd88}:		p = 14'd8360;
            {7'd95,7'd89}:		p = 14'd8455;
            {7'd95,7'd90}:		p = 14'd8550;
            {7'd95,7'd91}:		p = 14'd8645;
            {7'd95,7'd92}:		p = 14'd8740;
            {7'd95,7'd93}:		p = 14'd8835;
            {7'd95,7'd94}:		p = 14'd8930;
            {7'd95,7'd95}:		p = 14'd9025;
            {7'd95,7'd96}:		p = 14'd9120;
            {7'd95,7'd97}:		p = 14'd9215;
            {7'd95,7'd98}:		p = 14'd9310;
            {7'd95,7'd99}:		p = 14'd9405;
            {7'd95,7'd100}:		p = 14'd9500;
            {7'd95,7'd101}:		p = 14'd9595;
            {7'd95,7'd102}:		p = 14'd9690;
            {7'd95,7'd103}:		p = 14'd9785;
            {7'd95,7'd104}:		p = 14'd9880;
            {7'd95,7'd105}:		p = 14'd9975;
            {7'd95,7'd106}:		p = 14'd10070;
            {7'd95,7'd107}:		p = 14'd10165;
            {7'd95,7'd108}:		p = 14'd10260;
            {7'd95,7'd109}:		p = 14'd10355;
            {7'd95,7'd110}:		p = 14'd10450;
            {7'd95,7'd111}:		p = 14'd10545;
            {7'd95,7'd112}:		p = 14'd10640;
            {7'd95,7'd113}:		p = 14'd10735;
            {7'd95,7'd114}:		p = 14'd10830;
            {7'd95,7'd115}:		p = 14'd10925;
            {7'd95,7'd116}:		p = 14'd11020;
            {7'd95,7'd117}:		p = 14'd11115;
            {7'd95,7'd118}:		p = 14'd11210;
            {7'd95,7'd119}:		p = 14'd11305;
            {7'd95,7'd120}:		p = 14'd11400;
            {7'd95,7'd121}:		p = 14'd11495;
            {7'd95,7'd122}:		p = 14'd11590;
            {7'd95,7'd123}:		p = 14'd11685;
            {7'd95,7'd124}:		p = 14'd11780;
            {7'd95,7'd125}:		p = 14'd11875;
            {7'd95,7'd126}:		p = 14'd11970;
            {7'd95,7'd127}:		p = 14'd12065;
            {7'd96,7'd0}:		p = 14'd0;
            {7'd96,7'd1}:		p = 14'd96;
            {7'd96,7'd2}:		p = 14'd192;
            {7'd96,7'd3}:		p = 14'd288;
            {7'd96,7'd4}:		p = 14'd384;
            {7'd96,7'd5}:		p = 14'd480;
            {7'd96,7'd6}:		p = 14'd576;
            {7'd96,7'd7}:		p = 14'd672;
            {7'd96,7'd8}:		p = 14'd768;
            {7'd96,7'd9}:		p = 14'd864;
            {7'd96,7'd10}:		p = 14'd960;
            {7'd96,7'd11}:		p = 14'd1056;
            {7'd96,7'd12}:		p = 14'd1152;
            {7'd96,7'd13}:		p = 14'd1248;
            {7'd96,7'd14}:		p = 14'd1344;
            {7'd96,7'd15}:		p = 14'd1440;
            {7'd96,7'd16}:		p = 14'd1536;
            {7'd96,7'd17}:		p = 14'd1632;
            {7'd96,7'd18}:		p = 14'd1728;
            {7'd96,7'd19}:		p = 14'd1824;
            {7'd96,7'd20}:		p = 14'd1920;
            {7'd96,7'd21}:		p = 14'd2016;
            {7'd96,7'd22}:		p = 14'd2112;
            {7'd96,7'd23}:		p = 14'd2208;
            {7'd96,7'd24}:		p = 14'd2304;
            {7'd96,7'd25}:		p = 14'd2400;
            {7'd96,7'd26}:		p = 14'd2496;
            {7'd96,7'd27}:		p = 14'd2592;
            {7'd96,7'd28}:		p = 14'd2688;
            {7'd96,7'd29}:		p = 14'd2784;
            {7'd96,7'd30}:		p = 14'd2880;
            {7'd96,7'd31}:		p = 14'd2976;
            {7'd96,7'd32}:		p = 14'd3072;
            {7'd96,7'd33}:		p = 14'd3168;
            {7'd96,7'd34}:		p = 14'd3264;
            {7'd96,7'd35}:		p = 14'd3360;
            {7'd96,7'd36}:		p = 14'd3456;
            {7'd96,7'd37}:		p = 14'd3552;
            {7'd96,7'd38}:		p = 14'd3648;
            {7'd96,7'd39}:		p = 14'd3744;
            {7'd96,7'd40}:		p = 14'd3840;
            {7'd96,7'd41}:		p = 14'd3936;
            {7'd96,7'd42}:		p = 14'd4032;
            {7'd96,7'd43}:		p = 14'd4128;
            {7'd96,7'd44}:		p = 14'd4224;
            {7'd96,7'd45}:		p = 14'd4320;
            {7'd96,7'd46}:		p = 14'd4416;
            {7'd96,7'd47}:		p = 14'd4512;
            {7'd96,7'd48}:		p = 14'd4608;
            {7'd96,7'd49}:		p = 14'd4704;
            {7'd96,7'd50}:		p = 14'd4800;
            {7'd96,7'd51}:		p = 14'd4896;
            {7'd96,7'd52}:		p = 14'd4992;
            {7'd96,7'd53}:		p = 14'd5088;
            {7'd96,7'd54}:		p = 14'd5184;
            {7'd96,7'd55}:		p = 14'd5280;
            {7'd96,7'd56}:		p = 14'd5376;
            {7'd96,7'd57}:		p = 14'd5472;
            {7'd96,7'd58}:		p = 14'd5568;
            {7'd96,7'd59}:		p = 14'd5664;
            {7'd96,7'd60}:		p = 14'd5760;
            {7'd96,7'd61}:		p = 14'd5856;
            {7'd96,7'd62}:		p = 14'd5952;
            {7'd96,7'd63}:		p = 14'd6048;
            {7'd96,7'd64}:		p = 14'd6144;
            {7'd96,7'd65}:		p = 14'd6240;
            {7'd96,7'd66}:		p = 14'd6336;
            {7'd96,7'd67}:		p = 14'd6432;
            {7'd96,7'd68}:		p = 14'd6528;
            {7'd96,7'd69}:		p = 14'd6624;
            {7'd96,7'd70}:		p = 14'd6720;
            {7'd96,7'd71}:		p = 14'd6816;
            {7'd96,7'd72}:		p = 14'd6912;
            {7'd96,7'd73}:		p = 14'd7008;
            {7'd96,7'd74}:		p = 14'd7104;
            {7'd96,7'd75}:		p = 14'd7200;
            {7'd96,7'd76}:		p = 14'd7296;
            {7'd96,7'd77}:		p = 14'd7392;
            {7'd96,7'd78}:		p = 14'd7488;
            {7'd96,7'd79}:		p = 14'd7584;
            {7'd96,7'd80}:		p = 14'd7680;
            {7'd96,7'd81}:		p = 14'd7776;
            {7'd96,7'd82}:		p = 14'd7872;
            {7'd96,7'd83}:		p = 14'd7968;
            {7'd96,7'd84}:		p = 14'd8064;
            {7'd96,7'd85}:		p = 14'd8160;
            {7'd96,7'd86}:		p = 14'd8256;
            {7'd96,7'd87}:		p = 14'd8352;
            {7'd96,7'd88}:		p = 14'd8448;
            {7'd96,7'd89}:		p = 14'd8544;
            {7'd96,7'd90}:		p = 14'd8640;
            {7'd96,7'd91}:		p = 14'd8736;
            {7'd96,7'd92}:		p = 14'd8832;
            {7'd96,7'd93}:		p = 14'd8928;
            {7'd96,7'd94}:		p = 14'd9024;
            {7'd96,7'd95}:		p = 14'd9120;
            {7'd96,7'd96}:		p = 14'd9216;
            {7'd96,7'd97}:		p = 14'd9312;
            {7'd96,7'd98}:		p = 14'd9408;
            {7'd96,7'd99}:		p = 14'd9504;
            {7'd96,7'd100}:		p = 14'd9600;
            {7'd96,7'd101}:		p = 14'd9696;
            {7'd96,7'd102}:		p = 14'd9792;
            {7'd96,7'd103}:		p = 14'd9888;
            {7'd96,7'd104}:		p = 14'd9984;
            {7'd96,7'd105}:		p = 14'd10080;
            {7'd96,7'd106}:		p = 14'd10176;
            {7'd96,7'd107}:		p = 14'd10272;
            {7'd96,7'd108}:		p = 14'd10368;
            {7'd96,7'd109}:		p = 14'd10464;
            {7'd96,7'd110}:		p = 14'd10560;
            {7'd96,7'd111}:		p = 14'd10656;
            {7'd96,7'd112}:		p = 14'd10752;
            {7'd96,7'd113}:		p = 14'd10848;
            {7'd96,7'd114}:		p = 14'd10944;
            {7'd96,7'd115}:		p = 14'd11040;
            {7'd96,7'd116}:		p = 14'd11136;
            {7'd96,7'd117}:		p = 14'd11232;
            {7'd96,7'd118}:		p = 14'd11328;
            {7'd96,7'd119}:		p = 14'd11424;
            {7'd96,7'd120}:		p = 14'd11520;
            {7'd96,7'd121}:		p = 14'd11616;
            {7'd96,7'd122}:		p = 14'd11712;
            {7'd96,7'd123}:		p = 14'd11808;
            {7'd96,7'd124}:		p = 14'd11904;
            {7'd96,7'd125}:		p = 14'd12000;
            {7'd96,7'd126}:		p = 14'd12096;
            {7'd96,7'd127}:		p = 14'd12192;
            {7'd97,7'd0}:		p = 14'd0;
            {7'd97,7'd1}:		p = 14'd97;
            {7'd97,7'd2}:		p = 14'd194;
            {7'd97,7'd3}:		p = 14'd291;
            {7'd97,7'd4}:		p = 14'd388;
            {7'd97,7'd5}:		p = 14'd485;
            {7'd97,7'd6}:		p = 14'd582;
            {7'd97,7'd7}:		p = 14'd679;
            {7'd97,7'd8}:		p = 14'd776;
            {7'd97,7'd9}:		p = 14'd873;
            {7'd97,7'd10}:		p = 14'd970;
            {7'd97,7'd11}:		p = 14'd1067;
            {7'd97,7'd12}:		p = 14'd1164;
            {7'd97,7'd13}:		p = 14'd1261;
            {7'd97,7'd14}:		p = 14'd1358;
            {7'd97,7'd15}:		p = 14'd1455;
            {7'd97,7'd16}:		p = 14'd1552;
            {7'd97,7'd17}:		p = 14'd1649;
            {7'd97,7'd18}:		p = 14'd1746;
            {7'd97,7'd19}:		p = 14'd1843;
            {7'd97,7'd20}:		p = 14'd1940;
            {7'd97,7'd21}:		p = 14'd2037;
            {7'd97,7'd22}:		p = 14'd2134;
            {7'd97,7'd23}:		p = 14'd2231;
            {7'd97,7'd24}:		p = 14'd2328;
            {7'd97,7'd25}:		p = 14'd2425;
            {7'd97,7'd26}:		p = 14'd2522;
            {7'd97,7'd27}:		p = 14'd2619;
            {7'd97,7'd28}:		p = 14'd2716;
            {7'd97,7'd29}:		p = 14'd2813;
            {7'd97,7'd30}:		p = 14'd2910;
            {7'd97,7'd31}:		p = 14'd3007;
            {7'd97,7'd32}:		p = 14'd3104;
            {7'd97,7'd33}:		p = 14'd3201;
            {7'd97,7'd34}:		p = 14'd3298;
            {7'd97,7'd35}:		p = 14'd3395;
            {7'd97,7'd36}:		p = 14'd3492;
            {7'd97,7'd37}:		p = 14'd3589;
            {7'd97,7'd38}:		p = 14'd3686;
            {7'd97,7'd39}:		p = 14'd3783;
            {7'd97,7'd40}:		p = 14'd3880;
            {7'd97,7'd41}:		p = 14'd3977;
            {7'd97,7'd42}:		p = 14'd4074;
            {7'd97,7'd43}:		p = 14'd4171;
            {7'd97,7'd44}:		p = 14'd4268;
            {7'd97,7'd45}:		p = 14'd4365;
            {7'd97,7'd46}:		p = 14'd4462;
            {7'd97,7'd47}:		p = 14'd4559;
            {7'd97,7'd48}:		p = 14'd4656;
            {7'd97,7'd49}:		p = 14'd4753;
            {7'd97,7'd50}:		p = 14'd4850;
            {7'd97,7'd51}:		p = 14'd4947;
            {7'd97,7'd52}:		p = 14'd5044;
            {7'd97,7'd53}:		p = 14'd5141;
            {7'd97,7'd54}:		p = 14'd5238;
            {7'd97,7'd55}:		p = 14'd5335;
            {7'd97,7'd56}:		p = 14'd5432;
            {7'd97,7'd57}:		p = 14'd5529;
            {7'd97,7'd58}:		p = 14'd5626;
            {7'd97,7'd59}:		p = 14'd5723;
            {7'd97,7'd60}:		p = 14'd5820;
            {7'd97,7'd61}:		p = 14'd5917;
            {7'd97,7'd62}:		p = 14'd6014;
            {7'd97,7'd63}:		p = 14'd6111;
            {7'd97,7'd64}:		p = 14'd6208;
            {7'd97,7'd65}:		p = 14'd6305;
            {7'd97,7'd66}:		p = 14'd6402;
            {7'd97,7'd67}:		p = 14'd6499;
            {7'd97,7'd68}:		p = 14'd6596;
            {7'd97,7'd69}:		p = 14'd6693;
            {7'd97,7'd70}:		p = 14'd6790;
            {7'd97,7'd71}:		p = 14'd6887;
            {7'd97,7'd72}:		p = 14'd6984;
            {7'd97,7'd73}:		p = 14'd7081;
            {7'd97,7'd74}:		p = 14'd7178;
            {7'd97,7'd75}:		p = 14'd7275;
            {7'd97,7'd76}:		p = 14'd7372;
            {7'd97,7'd77}:		p = 14'd7469;
            {7'd97,7'd78}:		p = 14'd7566;
            {7'd97,7'd79}:		p = 14'd7663;
            {7'd97,7'd80}:		p = 14'd7760;
            {7'd97,7'd81}:		p = 14'd7857;
            {7'd97,7'd82}:		p = 14'd7954;
            {7'd97,7'd83}:		p = 14'd8051;
            {7'd97,7'd84}:		p = 14'd8148;
            {7'd97,7'd85}:		p = 14'd8245;
            {7'd97,7'd86}:		p = 14'd8342;
            {7'd97,7'd87}:		p = 14'd8439;
            {7'd97,7'd88}:		p = 14'd8536;
            {7'd97,7'd89}:		p = 14'd8633;
            {7'd97,7'd90}:		p = 14'd8730;
            {7'd97,7'd91}:		p = 14'd8827;
            {7'd97,7'd92}:		p = 14'd8924;
            {7'd97,7'd93}:		p = 14'd9021;
            {7'd97,7'd94}:		p = 14'd9118;
            {7'd97,7'd95}:		p = 14'd9215;
            {7'd97,7'd96}:		p = 14'd9312;
            {7'd97,7'd97}:		p = 14'd9409;
            {7'd97,7'd98}:		p = 14'd9506;
            {7'd97,7'd99}:		p = 14'd9603;
            {7'd97,7'd100}:		p = 14'd9700;
            {7'd97,7'd101}:		p = 14'd9797;
            {7'd97,7'd102}:		p = 14'd9894;
            {7'd97,7'd103}:		p = 14'd9991;
            {7'd97,7'd104}:		p = 14'd10088;
            {7'd97,7'd105}:		p = 14'd10185;
            {7'd97,7'd106}:		p = 14'd10282;
            {7'd97,7'd107}:		p = 14'd10379;
            {7'd97,7'd108}:		p = 14'd10476;
            {7'd97,7'd109}:		p = 14'd10573;
            {7'd97,7'd110}:		p = 14'd10670;
            {7'd97,7'd111}:		p = 14'd10767;
            {7'd97,7'd112}:		p = 14'd10864;
            {7'd97,7'd113}:		p = 14'd10961;
            {7'd97,7'd114}:		p = 14'd11058;
            {7'd97,7'd115}:		p = 14'd11155;
            {7'd97,7'd116}:		p = 14'd11252;
            {7'd97,7'd117}:		p = 14'd11349;
            {7'd97,7'd118}:		p = 14'd11446;
            {7'd97,7'd119}:		p = 14'd11543;
            {7'd97,7'd120}:		p = 14'd11640;
            {7'd97,7'd121}:		p = 14'd11737;
            {7'd97,7'd122}:		p = 14'd11834;
            {7'd97,7'd123}:		p = 14'd11931;
            {7'd97,7'd124}:		p = 14'd12028;
            {7'd97,7'd125}:		p = 14'd12125;
            {7'd97,7'd126}:		p = 14'd12222;
            {7'd97,7'd127}:		p = 14'd12319;
            {7'd98,7'd0}:		p = 14'd0;
            {7'd98,7'd1}:		p = 14'd98;
            {7'd98,7'd2}:		p = 14'd196;
            {7'd98,7'd3}:		p = 14'd294;
            {7'd98,7'd4}:		p = 14'd392;
            {7'd98,7'd5}:		p = 14'd490;
            {7'd98,7'd6}:		p = 14'd588;
            {7'd98,7'd7}:		p = 14'd686;
            {7'd98,7'd8}:		p = 14'd784;
            {7'd98,7'd9}:		p = 14'd882;
            {7'd98,7'd10}:		p = 14'd980;
            {7'd98,7'd11}:		p = 14'd1078;
            {7'd98,7'd12}:		p = 14'd1176;
            {7'd98,7'd13}:		p = 14'd1274;
            {7'd98,7'd14}:		p = 14'd1372;
            {7'd98,7'd15}:		p = 14'd1470;
            {7'd98,7'd16}:		p = 14'd1568;
            {7'd98,7'd17}:		p = 14'd1666;
            {7'd98,7'd18}:		p = 14'd1764;
            {7'd98,7'd19}:		p = 14'd1862;
            {7'd98,7'd20}:		p = 14'd1960;
            {7'd98,7'd21}:		p = 14'd2058;
            {7'd98,7'd22}:		p = 14'd2156;
            {7'd98,7'd23}:		p = 14'd2254;
            {7'd98,7'd24}:		p = 14'd2352;
            {7'd98,7'd25}:		p = 14'd2450;
            {7'd98,7'd26}:		p = 14'd2548;
            {7'd98,7'd27}:		p = 14'd2646;
            {7'd98,7'd28}:		p = 14'd2744;
            {7'd98,7'd29}:		p = 14'd2842;
            {7'd98,7'd30}:		p = 14'd2940;
            {7'd98,7'd31}:		p = 14'd3038;
            {7'd98,7'd32}:		p = 14'd3136;
            {7'd98,7'd33}:		p = 14'd3234;
            {7'd98,7'd34}:		p = 14'd3332;
            {7'd98,7'd35}:		p = 14'd3430;
            {7'd98,7'd36}:		p = 14'd3528;
            {7'd98,7'd37}:		p = 14'd3626;
            {7'd98,7'd38}:		p = 14'd3724;
            {7'd98,7'd39}:		p = 14'd3822;
            {7'd98,7'd40}:		p = 14'd3920;
            {7'd98,7'd41}:		p = 14'd4018;
            {7'd98,7'd42}:		p = 14'd4116;
            {7'd98,7'd43}:		p = 14'd4214;
            {7'd98,7'd44}:		p = 14'd4312;
            {7'd98,7'd45}:		p = 14'd4410;
            {7'd98,7'd46}:		p = 14'd4508;
            {7'd98,7'd47}:		p = 14'd4606;
            {7'd98,7'd48}:		p = 14'd4704;
            {7'd98,7'd49}:		p = 14'd4802;
            {7'd98,7'd50}:		p = 14'd4900;
            {7'd98,7'd51}:		p = 14'd4998;
            {7'd98,7'd52}:		p = 14'd5096;
            {7'd98,7'd53}:		p = 14'd5194;
            {7'd98,7'd54}:		p = 14'd5292;
            {7'd98,7'd55}:		p = 14'd5390;
            {7'd98,7'd56}:		p = 14'd5488;
            {7'd98,7'd57}:		p = 14'd5586;
            {7'd98,7'd58}:		p = 14'd5684;
            {7'd98,7'd59}:		p = 14'd5782;
            {7'd98,7'd60}:		p = 14'd5880;
            {7'd98,7'd61}:		p = 14'd5978;
            {7'd98,7'd62}:		p = 14'd6076;
            {7'd98,7'd63}:		p = 14'd6174;
            {7'd98,7'd64}:		p = 14'd6272;
            {7'd98,7'd65}:		p = 14'd6370;
            {7'd98,7'd66}:		p = 14'd6468;
            {7'd98,7'd67}:		p = 14'd6566;
            {7'd98,7'd68}:		p = 14'd6664;
            {7'd98,7'd69}:		p = 14'd6762;
            {7'd98,7'd70}:		p = 14'd6860;
            {7'd98,7'd71}:		p = 14'd6958;
            {7'd98,7'd72}:		p = 14'd7056;
            {7'd98,7'd73}:		p = 14'd7154;
            {7'd98,7'd74}:		p = 14'd7252;
            {7'd98,7'd75}:		p = 14'd7350;
            {7'd98,7'd76}:		p = 14'd7448;
            {7'd98,7'd77}:		p = 14'd7546;
            {7'd98,7'd78}:		p = 14'd7644;
            {7'd98,7'd79}:		p = 14'd7742;
            {7'd98,7'd80}:		p = 14'd7840;
            {7'd98,7'd81}:		p = 14'd7938;
            {7'd98,7'd82}:		p = 14'd8036;
            {7'd98,7'd83}:		p = 14'd8134;
            {7'd98,7'd84}:		p = 14'd8232;
            {7'd98,7'd85}:		p = 14'd8330;
            {7'd98,7'd86}:		p = 14'd8428;
            {7'd98,7'd87}:		p = 14'd8526;
            {7'd98,7'd88}:		p = 14'd8624;
            {7'd98,7'd89}:		p = 14'd8722;
            {7'd98,7'd90}:		p = 14'd8820;
            {7'd98,7'd91}:		p = 14'd8918;
            {7'd98,7'd92}:		p = 14'd9016;
            {7'd98,7'd93}:		p = 14'd9114;
            {7'd98,7'd94}:		p = 14'd9212;
            {7'd98,7'd95}:		p = 14'd9310;
            {7'd98,7'd96}:		p = 14'd9408;
            {7'd98,7'd97}:		p = 14'd9506;
            {7'd98,7'd98}:		p = 14'd9604;
            {7'd98,7'd99}:		p = 14'd9702;
            {7'd98,7'd100}:		p = 14'd9800;
            {7'd98,7'd101}:		p = 14'd9898;
            {7'd98,7'd102}:		p = 14'd9996;
            {7'd98,7'd103}:		p = 14'd10094;
            {7'd98,7'd104}:		p = 14'd10192;
            {7'd98,7'd105}:		p = 14'd10290;
            {7'd98,7'd106}:		p = 14'd10388;
            {7'd98,7'd107}:		p = 14'd10486;
            {7'd98,7'd108}:		p = 14'd10584;
            {7'd98,7'd109}:		p = 14'd10682;
            {7'd98,7'd110}:		p = 14'd10780;
            {7'd98,7'd111}:		p = 14'd10878;
            {7'd98,7'd112}:		p = 14'd10976;
            {7'd98,7'd113}:		p = 14'd11074;
            {7'd98,7'd114}:		p = 14'd11172;
            {7'd98,7'd115}:		p = 14'd11270;
            {7'd98,7'd116}:		p = 14'd11368;
            {7'd98,7'd117}:		p = 14'd11466;
            {7'd98,7'd118}:		p = 14'd11564;
            {7'd98,7'd119}:		p = 14'd11662;
            {7'd98,7'd120}:		p = 14'd11760;
            {7'd98,7'd121}:		p = 14'd11858;
            {7'd98,7'd122}:		p = 14'd11956;
            {7'd98,7'd123}:		p = 14'd12054;
            {7'd98,7'd124}:		p = 14'd12152;
            {7'd98,7'd125}:		p = 14'd12250;
            {7'd98,7'd126}:		p = 14'd12348;
            {7'd98,7'd127}:		p = 14'd12446;
            {7'd99,7'd0}:		p = 14'd0;
            {7'd99,7'd1}:		p = 14'd99;
            {7'd99,7'd2}:		p = 14'd198;
            {7'd99,7'd3}:		p = 14'd297;
            {7'd99,7'd4}:		p = 14'd396;
            {7'd99,7'd5}:		p = 14'd495;
            {7'd99,7'd6}:		p = 14'd594;
            {7'd99,7'd7}:		p = 14'd693;
            {7'd99,7'd8}:		p = 14'd792;
            {7'd99,7'd9}:		p = 14'd891;
            {7'd99,7'd10}:		p = 14'd990;
            {7'd99,7'd11}:		p = 14'd1089;
            {7'd99,7'd12}:		p = 14'd1188;
            {7'd99,7'd13}:		p = 14'd1287;
            {7'd99,7'd14}:		p = 14'd1386;
            {7'd99,7'd15}:		p = 14'd1485;
            {7'd99,7'd16}:		p = 14'd1584;
            {7'd99,7'd17}:		p = 14'd1683;
            {7'd99,7'd18}:		p = 14'd1782;
            {7'd99,7'd19}:		p = 14'd1881;
            {7'd99,7'd20}:		p = 14'd1980;
            {7'd99,7'd21}:		p = 14'd2079;
            {7'd99,7'd22}:		p = 14'd2178;
            {7'd99,7'd23}:		p = 14'd2277;
            {7'd99,7'd24}:		p = 14'd2376;
            {7'd99,7'd25}:		p = 14'd2475;
            {7'd99,7'd26}:		p = 14'd2574;
            {7'd99,7'd27}:		p = 14'd2673;
            {7'd99,7'd28}:		p = 14'd2772;
            {7'd99,7'd29}:		p = 14'd2871;
            {7'd99,7'd30}:		p = 14'd2970;
            {7'd99,7'd31}:		p = 14'd3069;
            {7'd99,7'd32}:		p = 14'd3168;
            {7'd99,7'd33}:		p = 14'd3267;
            {7'd99,7'd34}:		p = 14'd3366;
            {7'd99,7'd35}:		p = 14'd3465;
            {7'd99,7'd36}:		p = 14'd3564;
            {7'd99,7'd37}:		p = 14'd3663;
            {7'd99,7'd38}:		p = 14'd3762;
            {7'd99,7'd39}:		p = 14'd3861;
            {7'd99,7'd40}:		p = 14'd3960;
            {7'd99,7'd41}:		p = 14'd4059;
            {7'd99,7'd42}:		p = 14'd4158;
            {7'd99,7'd43}:		p = 14'd4257;
            {7'd99,7'd44}:		p = 14'd4356;
            {7'd99,7'd45}:		p = 14'd4455;
            {7'd99,7'd46}:		p = 14'd4554;
            {7'd99,7'd47}:		p = 14'd4653;
            {7'd99,7'd48}:		p = 14'd4752;
            {7'd99,7'd49}:		p = 14'd4851;
            {7'd99,7'd50}:		p = 14'd4950;
            {7'd99,7'd51}:		p = 14'd5049;
            {7'd99,7'd52}:		p = 14'd5148;
            {7'd99,7'd53}:		p = 14'd5247;
            {7'd99,7'd54}:		p = 14'd5346;
            {7'd99,7'd55}:		p = 14'd5445;
            {7'd99,7'd56}:		p = 14'd5544;
            {7'd99,7'd57}:		p = 14'd5643;
            {7'd99,7'd58}:		p = 14'd5742;
            {7'd99,7'd59}:		p = 14'd5841;
            {7'd99,7'd60}:		p = 14'd5940;
            {7'd99,7'd61}:		p = 14'd6039;
            {7'd99,7'd62}:		p = 14'd6138;
            {7'd99,7'd63}:		p = 14'd6237;
            {7'd99,7'd64}:		p = 14'd6336;
            {7'd99,7'd65}:		p = 14'd6435;
            {7'd99,7'd66}:		p = 14'd6534;
            {7'd99,7'd67}:		p = 14'd6633;
            {7'd99,7'd68}:		p = 14'd6732;
            {7'd99,7'd69}:		p = 14'd6831;
            {7'd99,7'd70}:		p = 14'd6930;
            {7'd99,7'd71}:		p = 14'd7029;
            {7'd99,7'd72}:		p = 14'd7128;
            {7'd99,7'd73}:		p = 14'd7227;
            {7'd99,7'd74}:		p = 14'd7326;
            {7'd99,7'd75}:		p = 14'd7425;
            {7'd99,7'd76}:		p = 14'd7524;
            {7'd99,7'd77}:		p = 14'd7623;
            {7'd99,7'd78}:		p = 14'd7722;
            {7'd99,7'd79}:		p = 14'd7821;
            {7'd99,7'd80}:		p = 14'd7920;
            {7'd99,7'd81}:		p = 14'd8019;
            {7'd99,7'd82}:		p = 14'd8118;
            {7'd99,7'd83}:		p = 14'd8217;
            {7'd99,7'd84}:		p = 14'd8316;
            {7'd99,7'd85}:		p = 14'd8415;
            {7'd99,7'd86}:		p = 14'd8514;
            {7'd99,7'd87}:		p = 14'd8613;
            {7'd99,7'd88}:		p = 14'd8712;
            {7'd99,7'd89}:		p = 14'd8811;
            {7'd99,7'd90}:		p = 14'd8910;
            {7'd99,7'd91}:		p = 14'd9009;
            {7'd99,7'd92}:		p = 14'd9108;
            {7'd99,7'd93}:		p = 14'd9207;
            {7'd99,7'd94}:		p = 14'd9306;
            {7'd99,7'd95}:		p = 14'd9405;
            {7'd99,7'd96}:		p = 14'd9504;
            {7'd99,7'd97}:		p = 14'd9603;
            {7'd99,7'd98}:		p = 14'd9702;
            {7'd99,7'd99}:		p = 14'd9801;
            {7'd99,7'd100}:		p = 14'd9900;
            {7'd99,7'd101}:		p = 14'd9999;
            {7'd99,7'd102}:		p = 14'd10098;
            {7'd99,7'd103}:		p = 14'd10197;
            {7'd99,7'd104}:		p = 14'd10296;
            {7'd99,7'd105}:		p = 14'd10395;
            {7'd99,7'd106}:		p = 14'd10494;
            {7'd99,7'd107}:		p = 14'd10593;
            {7'd99,7'd108}:		p = 14'd10692;
            {7'd99,7'd109}:		p = 14'd10791;
            {7'd99,7'd110}:		p = 14'd10890;
            {7'd99,7'd111}:		p = 14'd10989;
            {7'd99,7'd112}:		p = 14'd11088;
            {7'd99,7'd113}:		p = 14'd11187;
            {7'd99,7'd114}:		p = 14'd11286;
            {7'd99,7'd115}:		p = 14'd11385;
            {7'd99,7'd116}:		p = 14'd11484;
            {7'd99,7'd117}:		p = 14'd11583;
            {7'd99,7'd118}:		p = 14'd11682;
            {7'd99,7'd119}:		p = 14'd11781;
            {7'd99,7'd120}:		p = 14'd11880;
            {7'd99,7'd121}:		p = 14'd11979;
            {7'd99,7'd122}:		p = 14'd12078;
            {7'd99,7'd123}:		p = 14'd12177;
            {7'd99,7'd124}:		p = 14'd12276;
            {7'd99,7'd125}:		p = 14'd12375;
            {7'd99,7'd126}:		p = 14'd12474;
            {7'd99,7'd127}:		p = 14'd12573;
            {7'd100,7'd0}:		p = 14'd0;
            {7'd100,7'd1}:		p = 14'd100;
            {7'd100,7'd2}:		p = 14'd200;
            {7'd100,7'd3}:		p = 14'd300;
            {7'd100,7'd4}:		p = 14'd400;
            {7'd100,7'd5}:		p = 14'd500;
            {7'd100,7'd6}:		p = 14'd600;
            {7'd100,7'd7}:		p = 14'd700;
            {7'd100,7'd8}:		p = 14'd800;
            {7'd100,7'd9}:		p = 14'd900;
            {7'd100,7'd10}:		p = 14'd1000;
            {7'd100,7'd11}:		p = 14'd1100;
            {7'd100,7'd12}:		p = 14'd1200;
            {7'd100,7'd13}:		p = 14'd1300;
            {7'd100,7'd14}:		p = 14'd1400;
            {7'd100,7'd15}:		p = 14'd1500;
            {7'd100,7'd16}:		p = 14'd1600;
            {7'd100,7'd17}:		p = 14'd1700;
            {7'd100,7'd18}:		p = 14'd1800;
            {7'd100,7'd19}:		p = 14'd1900;
            {7'd100,7'd20}:		p = 14'd2000;
            {7'd100,7'd21}:		p = 14'd2100;
            {7'd100,7'd22}:		p = 14'd2200;
            {7'd100,7'd23}:		p = 14'd2300;
            {7'd100,7'd24}:		p = 14'd2400;
            {7'd100,7'd25}:		p = 14'd2500;
            {7'd100,7'd26}:		p = 14'd2600;
            {7'd100,7'd27}:		p = 14'd2700;
            {7'd100,7'd28}:		p = 14'd2800;
            {7'd100,7'd29}:		p = 14'd2900;
            {7'd100,7'd30}:		p = 14'd3000;
            {7'd100,7'd31}:		p = 14'd3100;
            {7'd100,7'd32}:		p = 14'd3200;
            {7'd100,7'd33}:		p = 14'd3300;
            {7'd100,7'd34}:		p = 14'd3400;
            {7'd100,7'd35}:		p = 14'd3500;
            {7'd100,7'd36}:		p = 14'd3600;
            {7'd100,7'd37}:		p = 14'd3700;
            {7'd100,7'd38}:		p = 14'd3800;
            {7'd100,7'd39}:		p = 14'd3900;
            {7'd100,7'd40}:		p = 14'd4000;
            {7'd100,7'd41}:		p = 14'd4100;
            {7'd100,7'd42}:		p = 14'd4200;
            {7'd100,7'd43}:		p = 14'd4300;
            {7'd100,7'd44}:		p = 14'd4400;
            {7'd100,7'd45}:		p = 14'd4500;
            {7'd100,7'd46}:		p = 14'd4600;
            {7'd100,7'd47}:		p = 14'd4700;
            {7'd100,7'd48}:		p = 14'd4800;
            {7'd100,7'd49}:		p = 14'd4900;
            {7'd100,7'd50}:		p = 14'd5000;
            {7'd100,7'd51}:		p = 14'd5100;
            {7'd100,7'd52}:		p = 14'd5200;
            {7'd100,7'd53}:		p = 14'd5300;
            {7'd100,7'd54}:		p = 14'd5400;
            {7'd100,7'd55}:		p = 14'd5500;
            {7'd100,7'd56}:		p = 14'd5600;
            {7'd100,7'd57}:		p = 14'd5700;
            {7'd100,7'd58}:		p = 14'd5800;
            {7'd100,7'd59}:		p = 14'd5900;
            {7'd100,7'd60}:		p = 14'd6000;
            {7'd100,7'd61}:		p = 14'd6100;
            {7'd100,7'd62}:		p = 14'd6200;
            {7'd100,7'd63}:		p = 14'd6300;
            {7'd100,7'd64}:		p = 14'd6400;
            {7'd100,7'd65}:		p = 14'd6500;
            {7'd100,7'd66}:		p = 14'd6600;
            {7'd100,7'd67}:		p = 14'd6700;
            {7'd100,7'd68}:		p = 14'd6800;
            {7'd100,7'd69}:		p = 14'd6900;
            {7'd100,7'd70}:		p = 14'd7000;
            {7'd100,7'd71}:		p = 14'd7100;
            {7'd100,7'd72}:		p = 14'd7200;
            {7'd100,7'd73}:		p = 14'd7300;
            {7'd100,7'd74}:		p = 14'd7400;
            {7'd100,7'd75}:		p = 14'd7500;
            {7'd100,7'd76}:		p = 14'd7600;
            {7'd100,7'd77}:		p = 14'd7700;
            {7'd100,7'd78}:		p = 14'd7800;
            {7'd100,7'd79}:		p = 14'd7900;
            {7'd100,7'd80}:		p = 14'd8000;
            {7'd100,7'd81}:		p = 14'd8100;
            {7'd100,7'd82}:		p = 14'd8200;
            {7'd100,7'd83}:		p = 14'd8300;
            {7'd100,7'd84}:		p = 14'd8400;
            {7'd100,7'd85}:		p = 14'd8500;
            {7'd100,7'd86}:		p = 14'd8600;
            {7'd100,7'd87}:		p = 14'd8700;
            {7'd100,7'd88}:		p = 14'd8800;
            {7'd100,7'd89}:		p = 14'd8900;
            {7'd100,7'd90}:		p = 14'd9000;
            {7'd100,7'd91}:		p = 14'd9100;
            {7'd100,7'd92}:		p = 14'd9200;
            {7'd100,7'd93}:		p = 14'd9300;
            {7'd100,7'd94}:		p = 14'd9400;
            {7'd100,7'd95}:		p = 14'd9500;
            {7'd100,7'd96}:		p = 14'd9600;
            {7'd100,7'd97}:		p = 14'd9700;
            {7'd100,7'd98}:		p = 14'd9800;
            {7'd100,7'd99}:		p = 14'd9900;
            {7'd100,7'd100}:		p = 14'd10000;
            {7'd100,7'd101}:		p = 14'd10100;
            {7'd100,7'd102}:		p = 14'd10200;
            {7'd100,7'd103}:		p = 14'd10300;
            {7'd100,7'd104}:		p = 14'd10400;
            {7'd100,7'd105}:		p = 14'd10500;
            {7'd100,7'd106}:		p = 14'd10600;
            {7'd100,7'd107}:		p = 14'd10700;
            {7'd100,7'd108}:		p = 14'd10800;
            {7'd100,7'd109}:		p = 14'd10900;
            {7'd100,7'd110}:		p = 14'd11000;
            {7'd100,7'd111}:		p = 14'd11100;
            {7'd100,7'd112}:		p = 14'd11200;
            {7'd100,7'd113}:		p = 14'd11300;
            {7'd100,7'd114}:		p = 14'd11400;
            {7'd100,7'd115}:		p = 14'd11500;
            {7'd100,7'd116}:		p = 14'd11600;
            {7'd100,7'd117}:		p = 14'd11700;
            {7'd100,7'd118}:		p = 14'd11800;
            {7'd100,7'd119}:		p = 14'd11900;
            {7'd100,7'd120}:		p = 14'd12000;
            {7'd100,7'd121}:		p = 14'd12100;
            {7'd100,7'd122}:		p = 14'd12200;
            {7'd100,7'd123}:		p = 14'd12300;
            {7'd100,7'd124}:		p = 14'd12400;
            {7'd100,7'd125}:		p = 14'd12500;
            {7'd100,7'd126}:		p = 14'd12600;
            {7'd100,7'd127}:		p = 14'd12700;
            {7'd101,7'd0}:		p = 14'd0;
            {7'd101,7'd1}:		p = 14'd101;
            {7'd101,7'd2}:		p = 14'd202;
            {7'd101,7'd3}:		p = 14'd303;
            {7'd101,7'd4}:		p = 14'd404;
            {7'd101,7'd5}:		p = 14'd505;
            {7'd101,7'd6}:		p = 14'd606;
            {7'd101,7'd7}:		p = 14'd707;
            {7'd101,7'd8}:		p = 14'd808;
            {7'd101,7'd9}:		p = 14'd909;
            {7'd101,7'd10}:		p = 14'd1010;
            {7'd101,7'd11}:		p = 14'd1111;
            {7'd101,7'd12}:		p = 14'd1212;
            {7'd101,7'd13}:		p = 14'd1313;
            {7'd101,7'd14}:		p = 14'd1414;
            {7'd101,7'd15}:		p = 14'd1515;
            {7'd101,7'd16}:		p = 14'd1616;
            {7'd101,7'd17}:		p = 14'd1717;
            {7'd101,7'd18}:		p = 14'd1818;
            {7'd101,7'd19}:		p = 14'd1919;
            {7'd101,7'd20}:		p = 14'd2020;
            {7'd101,7'd21}:		p = 14'd2121;
            {7'd101,7'd22}:		p = 14'd2222;
            {7'd101,7'd23}:		p = 14'd2323;
            {7'd101,7'd24}:		p = 14'd2424;
            {7'd101,7'd25}:		p = 14'd2525;
            {7'd101,7'd26}:		p = 14'd2626;
            {7'd101,7'd27}:		p = 14'd2727;
            {7'd101,7'd28}:		p = 14'd2828;
            {7'd101,7'd29}:		p = 14'd2929;
            {7'd101,7'd30}:		p = 14'd3030;
            {7'd101,7'd31}:		p = 14'd3131;
            {7'd101,7'd32}:		p = 14'd3232;
            {7'd101,7'd33}:		p = 14'd3333;
            {7'd101,7'd34}:		p = 14'd3434;
            {7'd101,7'd35}:		p = 14'd3535;
            {7'd101,7'd36}:		p = 14'd3636;
            {7'd101,7'd37}:		p = 14'd3737;
            {7'd101,7'd38}:		p = 14'd3838;
            {7'd101,7'd39}:		p = 14'd3939;
            {7'd101,7'd40}:		p = 14'd4040;
            {7'd101,7'd41}:		p = 14'd4141;
            {7'd101,7'd42}:		p = 14'd4242;
            {7'd101,7'd43}:		p = 14'd4343;
            {7'd101,7'd44}:		p = 14'd4444;
            {7'd101,7'd45}:		p = 14'd4545;
            {7'd101,7'd46}:		p = 14'd4646;
            {7'd101,7'd47}:		p = 14'd4747;
            {7'd101,7'd48}:		p = 14'd4848;
            {7'd101,7'd49}:		p = 14'd4949;
            {7'd101,7'd50}:		p = 14'd5050;
            {7'd101,7'd51}:		p = 14'd5151;
            {7'd101,7'd52}:		p = 14'd5252;
            {7'd101,7'd53}:		p = 14'd5353;
            {7'd101,7'd54}:		p = 14'd5454;
            {7'd101,7'd55}:		p = 14'd5555;
            {7'd101,7'd56}:		p = 14'd5656;
            {7'd101,7'd57}:		p = 14'd5757;
            {7'd101,7'd58}:		p = 14'd5858;
            {7'd101,7'd59}:		p = 14'd5959;
            {7'd101,7'd60}:		p = 14'd6060;
            {7'd101,7'd61}:		p = 14'd6161;
            {7'd101,7'd62}:		p = 14'd6262;
            {7'd101,7'd63}:		p = 14'd6363;
            {7'd101,7'd64}:		p = 14'd6464;
            {7'd101,7'd65}:		p = 14'd6565;
            {7'd101,7'd66}:		p = 14'd6666;
            {7'd101,7'd67}:		p = 14'd6767;
            {7'd101,7'd68}:		p = 14'd6868;
            {7'd101,7'd69}:		p = 14'd6969;
            {7'd101,7'd70}:		p = 14'd7070;
            {7'd101,7'd71}:		p = 14'd7171;
            {7'd101,7'd72}:		p = 14'd7272;
            {7'd101,7'd73}:		p = 14'd7373;
            {7'd101,7'd74}:		p = 14'd7474;
            {7'd101,7'd75}:		p = 14'd7575;
            {7'd101,7'd76}:		p = 14'd7676;
            {7'd101,7'd77}:		p = 14'd7777;
            {7'd101,7'd78}:		p = 14'd7878;
            {7'd101,7'd79}:		p = 14'd7979;
            {7'd101,7'd80}:		p = 14'd8080;
            {7'd101,7'd81}:		p = 14'd8181;
            {7'd101,7'd82}:		p = 14'd8282;
            {7'd101,7'd83}:		p = 14'd8383;
            {7'd101,7'd84}:		p = 14'd8484;
            {7'd101,7'd85}:		p = 14'd8585;
            {7'd101,7'd86}:		p = 14'd8686;
            {7'd101,7'd87}:		p = 14'd8787;
            {7'd101,7'd88}:		p = 14'd8888;
            {7'd101,7'd89}:		p = 14'd8989;
            {7'd101,7'd90}:		p = 14'd9090;
            {7'd101,7'd91}:		p = 14'd9191;
            {7'd101,7'd92}:		p = 14'd9292;
            {7'd101,7'd93}:		p = 14'd9393;
            {7'd101,7'd94}:		p = 14'd9494;
            {7'd101,7'd95}:		p = 14'd9595;
            {7'd101,7'd96}:		p = 14'd9696;
            {7'd101,7'd97}:		p = 14'd9797;
            {7'd101,7'd98}:		p = 14'd9898;
            {7'd101,7'd99}:		p = 14'd9999;
            {7'd101,7'd100}:		p = 14'd10100;
            {7'd101,7'd101}:		p = 14'd10201;
            {7'd101,7'd102}:		p = 14'd10302;
            {7'd101,7'd103}:		p = 14'd10403;
            {7'd101,7'd104}:		p = 14'd10504;
            {7'd101,7'd105}:		p = 14'd10605;
            {7'd101,7'd106}:		p = 14'd10706;
            {7'd101,7'd107}:		p = 14'd10807;
            {7'd101,7'd108}:		p = 14'd10908;
            {7'd101,7'd109}:		p = 14'd11009;
            {7'd101,7'd110}:		p = 14'd11110;
            {7'd101,7'd111}:		p = 14'd11211;
            {7'd101,7'd112}:		p = 14'd11312;
            {7'd101,7'd113}:		p = 14'd11413;
            {7'd101,7'd114}:		p = 14'd11514;
            {7'd101,7'd115}:		p = 14'd11615;
            {7'd101,7'd116}:		p = 14'd11716;
            {7'd101,7'd117}:		p = 14'd11817;
            {7'd101,7'd118}:		p = 14'd11918;
            {7'd101,7'd119}:		p = 14'd12019;
            {7'd101,7'd120}:		p = 14'd12120;
            {7'd101,7'd121}:		p = 14'd12221;
            {7'd101,7'd122}:		p = 14'd12322;
            {7'd101,7'd123}:		p = 14'd12423;
            {7'd101,7'd124}:		p = 14'd12524;
            {7'd101,7'd125}:		p = 14'd12625;
            {7'd101,7'd126}:		p = 14'd12726;
            {7'd101,7'd127}:		p = 14'd12827;
            {7'd102,7'd0}:		p = 14'd0;
            {7'd102,7'd1}:		p = 14'd102;
            {7'd102,7'd2}:		p = 14'd204;
            {7'd102,7'd3}:		p = 14'd306;
            {7'd102,7'd4}:		p = 14'd408;
            {7'd102,7'd5}:		p = 14'd510;
            {7'd102,7'd6}:		p = 14'd612;
            {7'd102,7'd7}:		p = 14'd714;
            {7'd102,7'd8}:		p = 14'd816;
            {7'd102,7'd9}:		p = 14'd918;
            {7'd102,7'd10}:		p = 14'd1020;
            {7'd102,7'd11}:		p = 14'd1122;
            {7'd102,7'd12}:		p = 14'd1224;
            {7'd102,7'd13}:		p = 14'd1326;
            {7'd102,7'd14}:		p = 14'd1428;
            {7'd102,7'd15}:		p = 14'd1530;
            {7'd102,7'd16}:		p = 14'd1632;
            {7'd102,7'd17}:		p = 14'd1734;
            {7'd102,7'd18}:		p = 14'd1836;
            {7'd102,7'd19}:		p = 14'd1938;
            {7'd102,7'd20}:		p = 14'd2040;
            {7'd102,7'd21}:		p = 14'd2142;
            {7'd102,7'd22}:		p = 14'd2244;
            {7'd102,7'd23}:		p = 14'd2346;
            {7'd102,7'd24}:		p = 14'd2448;
            {7'd102,7'd25}:		p = 14'd2550;
            {7'd102,7'd26}:		p = 14'd2652;
            {7'd102,7'd27}:		p = 14'd2754;
            {7'd102,7'd28}:		p = 14'd2856;
            {7'd102,7'd29}:		p = 14'd2958;
            {7'd102,7'd30}:		p = 14'd3060;
            {7'd102,7'd31}:		p = 14'd3162;
            {7'd102,7'd32}:		p = 14'd3264;
            {7'd102,7'd33}:		p = 14'd3366;
            {7'd102,7'd34}:		p = 14'd3468;
            {7'd102,7'd35}:		p = 14'd3570;
            {7'd102,7'd36}:		p = 14'd3672;
            {7'd102,7'd37}:		p = 14'd3774;
            {7'd102,7'd38}:		p = 14'd3876;
            {7'd102,7'd39}:		p = 14'd3978;
            {7'd102,7'd40}:		p = 14'd4080;
            {7'd102,7'd41}:		p = 14'd4182;
            {7'd102,7'd42}:		p = 14'd4284;
            {7'd102,7'd43}:		p = 14'd4386;
            {7'd102,7'd44}:		p = 14'd4488;
            {7'd102,7'd45}:		p = 14'd4590;
            {7'd102,7'd46}:		p = 14'd4692;
            {7'd102,7'd47}:		p = 14'd4794;
            {7'd102,7'd48}:		p = 14'd4896;
            {7'd102,7'd49}:		p = 14'd4998;
            {7'd102,7'd50}:		p = 14'd5100;
            {7'd102,7'd51}:		p = 14'd5202;
            {7'd102,7'd52}:		p = 14'd5304;
            {7'd102,7'd53}:		p = 14'd5406;
            {7'd102,7'd54}:		p = 14'd5508;
            {7'd102,7'd55}:		p = 14'd5610;
            {7'd102,7'd56}:		p = 14'd5712;
            {7'd102,7'd57}:		p = 14'd5814;
            {7'd102,7'd58}:		p = 14'd5916;
            {7'd102,7'd59}:		p = 14'd6018;
            {7'd102,7'd60}:		p = 14'd6120;
            {7'd102,7'd61}:		p = 14'd6222;
            {7'd102,7'd62}:		p = 14'd6324;
            {7'd102,7'd63}:		p = 14'd6426;
            {7'd102,7'd64}:		p = 14'd6528;
            {7'd102,7'd65}:		p = 14'd6630;
            {7'd102,7'd66}:		p = 14'd6732;
            {7'd102,7'd67}:		p = 14'd6834;
            {7'd102,7'd68}:		p = 14'd6936;
            {7'd102,7'd69}:		p = 14'd7038;
            {7'd102,7'd70}:		p = 14'd7140;
            {7'd102,7'd71}:		p = 14'd7242;
            {7'd102,7'd72}:		p = 14'd7344;
            {7'd102,7'd73}:		p = 14'd7446;
            {7'd102,7'd74}:		p = 14'd7548;
            {7'd102,7'd75}:		p = 14'd7650;
            {7'd102,7'd76}:		p = 14'd7752;
            {7'd102,7'd77}:		p = 14'd7854;
            {7'd102,7'd78}:		p = 14'd7956;
            {7'd102,7'd79}:		p = 14'd8058;
            {7'd102,7'd80}:		p = 14'd8160;
            {7'd102,7'd81}:		p = 14'd8262;
            {7'd102,7'd82}:		p = 14'd8364;
            {7'd102,7'd83}:		p = 14'd8466;
            {7'd102,7'd84}:		p = 14'd8568;
            {7'd102,7'd85}:		p = 14'd8670;
            {7'd102,7'd86}:		p = 14'd8772;
            {7'd102,7'd87}:		p = 14'd8874;
            {7'd102,7'd88}:		p = 14'd8976;
            {7'd102,7'd89}:		p = 14'd9078;
            {7'd102,7'd90}:		p = 14'd9180;
            {7'd102,7'd91}:		p = 14'd9282;
            {7'd102,7'd92}:		p = 14'd9384;
            {7'd102,7'd93}:		p = 14'd9486;
            {7'd102,7'd94}:		p = 14'd9588;
            {7'd102,7'd95}:		p = 14'd9690;
            {7'd102,7'd96}:		p = 14'd9792;
            {7'd102,7'd97}:		p = 14'd9894;
            {7'd102,7'd98}:		p = 14'd9996;
            {7'd102,7'd99}:		p = 14'd10098;
            {7'd102,7'd100}:		p = 14'd10200;
            {7'd102,7'd101}:		p = 14'd10302;
            {7'd102,7'd102}:		p = 14'd10404;
            {7'd102,7'd103}:		p = 14'd10506;
            {7'd102,7'd104}:		p = 14'd10608;
            {7'd102,7'd105}:		p = 14'd10710;
            {7'd102,7'd106}:		p = 14'd10812;
            {7'd102,7'd107}:		p = 14'd10914;
            {7'd102,7'd108}:		p = 14'd11016;
            {7'd102,7'd109}:		p = 14'd11118;
            {7'd102,7'd110}:		p = 14'd11220;
            {7'd102,7'd111}:		p = 14'd11322;
            {7'd102,7'd112}:		p = 14'd11424;
            {7'd102,7'd113}:		p = 14'd11526;
            {7'd102,7'd114}:		p = 14'd11628;
            {7'd102,7'd115}:		p = 14'd11730;
            {7'd102,7'd116}:		p = 14'd11832;
            {7'd102,7'd117}:		p = 14'd11934;
            {7'd102,7'd118}:		p = 14'd12036;
            {7'd102,7'd119}:		p = 14'd12138;
            {7'd102,7'd120}:		p = 14'd12240;
            {7'd102,7'd121}:		p = 14'd12342;
            {7'd102,7'd122}:		p = 14'd12444;
            {7'd102,7'd123}:		p = 14'd12546;
            {7'd102,7'd124}:		p = 14'd12648;
            {7'd102,7'd125}:		p = 14'd12750;
            {7'd102,7'd126}:		p = 14'd12852;
            {7'd102,7'd127}:		p = 14'd12954;
            {7'd103,7'd0}:		p = 14'd0;
            {7'd103,7'd1}:		p = 14'd103;
            {7'd103,7'd2}:		p = 14'd206;
            {7'd103,7'd3}:		p = 14'd309;
            {7'd103,7'd4}:		p = 14'd412;
            {7'd103,7'd5}:		p = 14'd515;
            {7'd103,7'd6}:		p = 14'd618;
            {7'd103,7'd7}:		p = 14'd721;
            {7'd103,7'd8}:		p = 14'd824;
            {7'd103,7'd9}:		p = 14'd927;
            {7'd103,7'd10}:		p = 14'd1030;
            {7'd103,7'd11}:		p = 14'd1133;
            {7'd103,7'd12}:		p = 14'd1236;
            {7'd103,7'd13}:		p = 14'd1339;
            {7'd103,7'd14}:		p = 14'd1442;
            {7'd103,7'd15}:		p = 14'd1545;
            {7'd103,7'd16}:		p = 14'd1648;
            {7'd103,7'd17}:		p = 14'd1751;
            {7'd103,7'd18}:		p = 14'd1854;
            {7'd103,7'd19}:		p = 14'd1957;
            {7'd103,7'd20}:		p = 14'd2060;
            {7'd103,7'd21}:		p = 14'd2163;
            {7'd103,7'd22}:		p = 14'd2266;
            {7'd103,7'd23}:		p = 14'd2369;
            {7'd103,7'd24}:		p = 14'd2472;
            {7'd103,7'd25}:		p = 14'd2575;
            {7'd103,7'd26}:		p = 14'd2678;
            {7'd103,7'd27}:		p = 14'd2781;
            {7'd103,7'd28}:		p = 14'd2884;
            {7'd103,7'd29}:		p = 14'd2987;
            {7'd103,7'd30}:		p = 14'd3090;
            {7'd103,7'd31}:		p = 14'd3193;
            {7'd103,7'd32}:		p = 14'd3296;
            {7'd103,7'd33}:		p = 14'd3399;
            {7'd103,7'd34}:		p = 14'd3502;
            {7'd103,7'd35}:		p = 14'd3605;
            {7'd103,7'd36}:		p = 14'd3708;
            {7'd103,7'd37}:		p = 14'd3811;
            {7'd103,7'd38}:		p = 14'd3914;
            {7'd103,7'd39}:		p = 14'd4017;
            {7'd103,7'd40}:		p = 14'd4120;
            {7'd103,7'd41}:		p = 14'd4223;
            {7'd103,7'd42}:		p = 14'd4326;
            {7'd103,7'd43}:		p = 14'd4429;
            {7'd103,7'd44}:		p = 14'd4532;
            {7'd103,7'd45}:		p = 14'd4635;
            {7'd103,7'd46}:		p = 14'd4738;
            {7'd103,7'd47}:		p = 14'd4841;
            {7'd103,7'd48}:		p = 14'd4944;
            {7'd103,7'd49}:		p = 14'd5047;
            {7'd103,7'd50}:		p = 14'd5150;
            {7'd103,7'd51}:		p = 14'd5253;
            {7'd103,7'd52}:		p = 14'd5356;
            {7'd103,7'd53}:		p = 14'd5459;
            {7'd103,7'd54}:		p = 14'd5562;
            {7'd103,7'd55}:		p = 14'd5665;
            {7'd103,7'd56}:		p = 14'd5768;
            {7'd103,7'd57}:		p = 14'd5871;
            {7'd103,7'd58}:		p = 14'd5974;
            {7'd103,7'd59}:		p = 14'd6077;
            {7'd103,7'd60}:		p = 14'd6180;
            {7'd103,7'd61}:		p = 14'd6283;
            {7'd103,7'd62}:		p = 14'd6386;
            {7'd103,7'd63}:		p = 14'd6489;
            {7'd103,7'd64}:		p = 14'd6592;
            {7'd103,7'd65}:		p = 14'd6695;
            {7'd103,7'd66}:		p = 14'd6798;
            {7'd103,7'd67}:		p = 14'd6901;
            {7'd103,7'd68}:		p = 14'd7004;
            {7'd103,7'd69}:		p = 14'd7107;
            {7'd103,7'd70}:		p = 14'd7210;
            {7'd103,7'd71}:		p = 14'd7313;
            {7'd103,7'd72}:		p = 14'd7416;
            {7'd103,7'd73}:		p = 14'd7519;
            {7'd103,7'd74}:		p = 14'd7622;
            {7'd103,7'd75}:		p = 14'd7725;
            {7'd103,7'd76}:		p = 14'd7828;
            {7'd103,7'd77}:		p = 14'd7931;
            {7'd103,7'd78}:		p = 14'd8034;
            {7'd103,7'd79}:		p = 14'd8137;
            {7'd103,7'd80}:		p = 14'd8240;
            {7'd103,7'd81}:		p = 14'd8343;
            {7'd103,7'd82}:		p = 14'd8446;
            {7'd103,7'd83}:		p = 14'd8549;
            {7'd103,7'd84}:		p = 14'd8652;
            {7'd103,7'd85}:		p = 14'd8755;
            {7'd103,7'd86}:		p = 14'd8858;
            {7'd103,7'd87}:		p = 14'd8961;
            {7'd103,7'd88}:		p = 14'd9064;
            {7'd103,7'd89}:		p = 14'd9167;
            {7'd103,7'd90}:		p = 14'd9270;
            {7'd103,7'd91}:		p = 14'd9373;
            {7'd103,7'd92}:		p = 14'd9476;
            {7'd103,7'd93}:		p = 14'd9579;
            {7'd103,7'd94}:		p = 14'd9682;
            {7'd103,7'd95}:		p = 14'd9785;
            {7'd103,7'd96}:		p = 14'd9888;
            {7'd103,7'd97}:		p = 14'd9991;
            {7'd103,7'd98}:		p = 14'd10094;
            {7'd103,7'd99}:		p = 14'd10197;
            {7'd103,7'd100}:		p = 14'd10300;
            {7'd103,7'd101}:		p = 14'd10403;
            {7'd103,7'd102}:		p = 14'd10506;
            {7'd103,7'd103}:		p = 14'd10609;
            {7'd103,7'd104}:		p = 14'd10712;
            {7'd103,7'd105}:		p = 14'd10815;
            {7'd103,7'd106}:		p = 14'd10918;
            {7'd103,7'd107}:		p = 14'd11021;
            {7'd103,7'd108}:		p = 14'd11124;
            {7'd103,7'd109}:		p = 14'd11227;
            {7'd103,7'd110}:		p = 14'd11330;
            {7'd103,7'd111}:		p = 14'd11433;
            {7'd103,7'd112}:		p = 14'd11536;
            {7'd103,7'd113}:		p = 14'd11639;
            {7'd103,7'd114}:		p = 14'd11742;
            {7'd103,7'd115}:		p = 14'd11845;
            {7'd103,7'd116}:		p = 14'd11948;
            {7'd103,7'd117}:		p = 14'd12051;
            {7'd103,7'd118}:		p = 14'd12154;
            {7'd103,7'd119}:		p = 14'd12257;
            {7'd103,7'd120}:		p = 14'd12360;
            {7'd103,7'd121}:		p = 14'd12463;
            {7'd103,7'd122}:		p = 14'd12566;
            {7'd103,7'd123}:		p = 14'd12669;
            {7'd103,7'd124}:		p = 14'd12772;
            {7'd103,7'd125}:		p = 14'd12875;
            {7'd103,7'd126}:		p = 14'd12978;
            {7'd103,7'd127}:		p = 14'd13081;
            {7'd104,7'd0}:		p = 14'd0;
            {7'd104,7'd1}:		p = 14'd104;
            {7'd104,7'd2}:		p = 14'd208;
            {7'd104,7'd3}:		p = 14'd312;
            {7'd104,7'd4}:		p = 14'd416;
            {7'd104,7'd5}:		p = 14'd520;
            {7'd104,7'd6}:		p = 14'd624;
            {7'd104,7'd7}:		p = 14'd728;
            {7'd104,7'd8}:		p = 14'd832;
            {7'd104,7'd9}:		p = 14'd936;
            {7'd104,7'd10}:		p = 14'd1040;
            {7'd104,7'd11}:		p = 14'd1144;
            {7'd104,7'd12}:		p = 14'd1248;
            {7'd104,7'd13}:		p = 14'd1352;
            {7'd104,7'd14}:		p = 14'd1456;
            {7'd104,7'd15}:		p = 14'd1560;
            {7'd104,7'd16}:		p = 14'd1664;
            {7'd104,7'd17}:		p = 14'd1768;
            {7'd104,7'd18}:		p = 14'd1872;
            {7'd104,7'd19}:		p = 14'd1976;
            {7'd104,7'd20}:		p = 14'd2080;
            {7'd104,7'd21}:		p = 14'd2184;
            {7'd104,7'd22}:		p = 14'd2288;
            {7'd104,7'd23}:		p = 14'd2392;
            {7'd104,7'd24}:		p = 14'd2496;
            {7'd104,7'd25}:		p = 14'd2600;
            {7'd104,7'd26}:		p = 14'd2704;
            {7'd104,7'd27}:		p = 14'd2808;
            {7'd104,7'd28}:		p = 14'd2912;
            {7'd104,7'd29}:		p = 14'd3016;
            {7'd104,7'd30}:		p = 14'd3120;
            {7'd104,7'd31}:		p = 14'd3224;
            {7'd104,7'd32}:		p = 14'd3328;
            {7'd104,7'd33}:		p = 14'd3432;
            {7'd104,7'd34}:		p = 14'd3536;
            {7'd104,7'd35}:		p = 14'd3640;
            {7'd104,7'd36}:		p = 14'd3744;
            {7'd104,7'd37}:		p = 14'd3848;
            {7'd104,7'd38}:		p = 14'd3952;
            {7'd104,7'd39}:		p = 14'd4056;
            {7'd104,7'd40}:		p = 14'd4160;
            {7'd104,7'd41}:		p = 14'd4264;
            {7'd104,7'd42}:		p = 14'd4368;
            {7'd104,7'd43}:		p = 14'd4472;
            {7'd104,7'd44}:		p = 14'd4576;
            {7'd104,7'd45}:		p = 14'd4680;
            {7'd104,7'd46}:		p = 14'd4784;
            {7'd104,7'd47}:		p = 14'd4888;
            {7'd104,7'd48}:		p = 14'd4992;
            {7'd104,7'd49}:		p = 14'd5096;
            {7'd104,7'd50}:		p = 14'd5200;
            {7'd104,7'd51}:		p = 14'd5304;
            {7'd104,7'd52}:		p = 14'd5408;
            {7'd104,7'd53}:		p = 14'd5512;
            {7'd104,7'd54}:		p = 14'd5616;
            {7'd104,7'd55}:		p = 14'd5720;
            {7'd104,7'd56}:		p = 14'd5824;
            {7'd104,7'd57}:		p = 14'd5928;
            {7'd104,7'd58}:		p = 14'd6032;
            {7'd104,7'd59}:		p = 14'd6136;
            {7'd104,7'd60}:		p = 14'd6240;
            {7'd104,7'd61}:		p = 14'd6344;
            {7'd104,7'd62}:		p = 14'd6448;
            {7'd104,7'd63}:		p = 14'd6552;
            {7'd104,7'd64}:		p = 14'd6656;
            {7'd104,7'd65}:		p = 14'd6760;
            {7'd104,7'd66}:		p = 14'd6864;
            {7'd104,7'd67}:		p = 14'd6968;
            {7'd104,7'd68}:		p = 14'd7072;
            {7'd104,7'd69}:		p = 14'd7176;
            {7'd104,7'd70}:		p = 14'd7280;
            {7'd104,7'd71}:		p = 14'd7384;
            {7'd104,7'd72}:		p = 14'd7488;
            {7'd104,7'd73}:		p = 14'd7592;
            {7'd104,7'd74}:		p = 14'd7696;
            {7'd104,7'd75}:		p = 14'd7800;
            {7'd104,7'd76}:		p = 14'd7904;
            {7'd104,7'd77}:		p = 14'd8008;
            {7'd104,7'd78}:		p = 14'd8112;
            {7'd104,7'd79}:		p = 14'd8216;
            {7'd104,7'd80}:		p = 14'd8320;
            {7'd104,7'd81}:		p = 14'd8424;
            {7'd104,7'd82}:		p = 14'd8528;
            {7'd104,7'd83}:		p = 14'd8632;
            {7'd104,7'd84}:		p = 14'd8736;
            {7'd104,7'd85}:		p = 14'd8840;
            {7'd104,7'd86}:		p = 14'd8944;
            {7'd104,7'd87}:		p = 14'd9048;
            {7'd104,7'd88}:		p = 14'd9152;
            {7'd104,7'd89}:		p = 14'd9256;
            {7'd104,7'd90}:		p = 14'd9360;
            {7'd104,7'd91}:		p = 14'd9464;
            {7'd104,7'd92}:		p = 14'd9568;
            {7'd104,7'd93}:		p = 14'd9672;
            {7'd104,7'd94}:		p = 14'd9776;
            {7'd104,7'd95}:		p = 14'd9880;
            {7'd104,7'd96}:		p = 14'd9984;
            {7'd104,7'd97}:		p = 14'd10088;
            {7'd104,7'd98}:		p = 14'd10192;
            {7'd104,7'd99}:		p = 14'd10296;
            {7'd104,7'd100}:		p = 14'd10400;
            {7'd104,7'd101}:		p = 14'd10504;
            {7'd104,7'd102}:		p = 14'd10608;
            {7'd104,7'd103}:		p = 14'd10712;
            {7'd104,7'd104}:		p = 14'd10816;
            {7'd104,7'd105}:		p = 14'd10920;
            {7'd104,7'd106}:		p = 14'd11024;
            {7'd104,7'd107}:		p = 14'd11128;
            {7'd104,7'd108}:		p = 14'd11232;
            {7'd104,7'd109}:		p = 14'd11336;
            {7'd104,7'd110}:		p = 14'd11440;
            {7'd104,7'd111}:		p = 14'd11544;
            {7'd104,7'd112}:		p = 14'd11648;
            {7'd104,7'd113}:		p = 14'd11752;
            {7'd104,7'd114}:		p = 14'd11856;
            {7'd104,7'd115}:		p = 14'd11960;
            {7'd104,7'd116}:		p = 14'd12064;
            {7'd104,7'd117}:		p = 14'd12168;
            {7'd104,7'd118}:		p = 14'd12272;
            {7'd104,7'd119}:		p = 14'd12376;
            {7'd104,7'd120}:		p = 14'd12480;
            {7'd104,7'd121}:		p = 14'd12584;
            {7'd104,7'd122}:		p = 14'd12688;
            {7'd104,7'd123}:		p = 14'd12792;
            {7'd104,7'd124}:		p = 14'd12896;
            {7'd104,7'd125}:		p = 14'd13000;
            {7'd104,7'd126}:		p = 14'd13104;
            {7'd104,7'd127}:		p = 14'd13208;
            {7'd105,7'd0}:		p = 14'd0;
            {7'd105,7'd1}:		p = 14'd105;
            {7'd105,7'd2}:		p = 14'd210;
            {7'd105,7'd3}:		p = 14'd315;
            {7'd105,7'd4}:		p = 14'd420;
            {7'd105,7'd5}:		p = 14'd525;
            {7'd105,7'd6}:		p = 14'd630;
            {7'd105,7'd7}:		p = 14'd735;
            {7'd105,7'd8}:		p = 14'd840;
            {7'd105,7'd9}:		p = 14'd945;
            {7'd105,7'd10}:		p = 14'd1050;
            {7'd105,7'd11}:		p = 14'd1155;
            {7'd105,7'd12}:		p = 14'd1260;
            {7'd105,7'd13}:		p = 14'd1365;
            {7'd105,7'd14}:		p = 14'd1470;
            {7'd105,7'd15}:		p = 14'd1575;
            {7'd105,7'd16}:		p = 14'd1680;
            {7'd105,7'd17}:		p = 14'd1785;
            {7'd105,7'd18}:		p = 14'd1890;
            {7'd105,7'd19}:		p = 14'd1995;
            {7'd105,7'd20}:		p = 14'd2100;
            {7'd105,7'd21}:		p = 14'd2205;
            {7'd105,7'd22}:		p = 14'd2310;
            {7'd105,7'd23}:		p = 14'd2415;
            {7'd105,7'd24}:		p = 14'd2520;
            {7'd105,7'd25}:		p = 14'd2625;
            {7'd105,7'd26}:		p = 14'd2730;
            {7'd105,7'd27}:		p = 14'd2835;
            {7'd105,7'd28}:		p = 14'd2940;
            {7'd105,7'd29}:		p = 14'd3045;
            {7'd105,7'd30}:		p = 14'd3150;
            {7'd105,7'd31}:		p = 14'd3255;
            {7'd105,7'd32}:		p = 14'd3360;
            {7'd105,7'd33}:		p = 14'd3465;
            {7'd105,7'd34}:		p = 14'd3570;
            {7'd105,7'd35}:		p = 14'd3675;
            {7'd105,7'd36}:		p = 14'd3780;
            {7'd105,7'd37}:		p = 14'd3885;
            {7'd105,7'd38}:		p = 14'd3990;
            {7'd105,7'd39}:		p = 14'd4095;
            {7'd105,7'd40}:		p = 14'd4200;
            {7'd105,7'd41}:		p = 14'd4305;
            {7'd105,7'd42}:		p = 14'd4410;
            {7'd105,7'd43}:		p = 14'd4515;
            {7'd105,7'd44}:		p = 14'd4620;
            {7'd105,7'd45}:		p = 14'd4725;
            {7'd105,7'd46}:		p = 14'd4830;
            {7'd105,7'd47}:		p = 14'd4935;
            {7'd105,7'd48}:		p = 14'd5040;
            {7'd105,7'd49}:		p = 14'd5145;
            {7'd105,7'd50}:		p = 14'd5250;
            {7'd105,7'd51}:		p = 14'd5355;
            {7'd105,7'd52}:		p = 14'd5460;
            {7'd105,7'd53}:		p = 14'd5565;
            {7'd105,7'd54}:		p = 14'd5670;
            {7'd105,7'd55}:		p = 14'd5775;
            {7'd105,7'd56}:		p = 14'd5880;
            {7'd105,7'd57}:		p = 14'd5985;
            {7'd105,7'd58}:		p = 14'd6090;
            {7'd105,7'd59}:		p = 14'd6195;
            {7'd105,7'd60}:		p = 14'd6300;
            {7'd105,7'd61}:		p = 14'd6405;
            {7'd105,7'd62}:		p = 14'd6510;
            {7'd105,7'd63}:		p = 14'd6615;
            {7'd105,7'd64}:		p = 14'd6720;
            {7'd105,7'd65}:		p = 14'd6825;
            {7'd105,7'd66}:		p = 14'd6930;
            {7'd105,7'd67}:		p = 14'd7035;
            {7'd105,7'd68}:		p = 14'd7140;
            {7'd105,7'd69}:		p = 14'd7245;
            {7'd105,7'd70}:		p = 14'd7350;
            {7'd105,7'd71}:		p = 14'd7455;
            {7'd105,7'd72}:		p = 14'd7560;
            {7'd105,7'd73}:		p = 14'd7665;
            {7'd105,7'd74}:		p = 14'd7770;
            {7'd105,7'd75}:		p = 14'd7875;
            {7'd105,7'd76}:		p = 14'd7980;
            {7'd105,7'd77}:		p = 14'd8085;
            {7'd105,7'd78}:		p = 14'd8190;
            {7'd105,7'd79}:		p = 14'd8295;
            {7'd105,7'd80}:		p = 14'd8400;
            {7'd105,7'd81}:		p = 14'd8505;
            {7'd105,7'd82}:		p = 14'd8610;
            {7'd105,7'd83}:		p = 14'd8715;
            {7'd105,7'd84}:		p = 14'd8820;
            {7'd105,7'd85}:		p = 14'd8925;
            {7'd105,7'd86}:		p = 14'd9030;
            {7'd105,7'd87}:		p = 14'd9135;
            {7'd105,7'd88}:		p = 14'd9240;
            {7'd105,7'd89}:		p = 14'd9345;
            {7'd105,7'd90}:		p = 14'd9450;
            {7'd105,7'd91}:		p = 14'd9555;
            {7'd105,7'd92}:		p = 14'd9660;
            {7'd105,7'd93}:		p = 14'd9765;
            {7'd105,7'd94}:		p = 14'd9870;
            {7'd105,7'd95}:		p = 14'd9975;
            {7'd105,7'd96}:		p = 14'd10080;
            {7'd105,7'd97}:		p = 14'd10185;
            {7'd105,7'd98}:		p = 14'd10290;
            {7'd105,7'd99}:		p = 14'd10395;
            {7'd105,7'd100}:		p = 14'd10500;
            {7'd105,7'd101}:		p = 14'd10605;
            {7'd105,7'd102}:		p = 14'd10710;
            {7'd105,7'd103}:		p = 14'd10815;
            {7'd105,7'd104}:		p = 14'd10920;
            {7'd105,7'd105}:		p = 14'd11025;
            {7'd105,7'd106}:		p = 14'd11130;
            {7'd105,7'd107}:		p = 14'd11235;
            {7'd105,7'd108}:		p = 14'd11340;
            {7'd105,7'd109}:		p = 14'd11445;
            {7'd105,7'd110}:		p = 14'd11550;
            {7'd105,7'd111}:		p = 14'd11655;
            {7'd105,7'd112}:		p = 14'd11760;
            {7'd105,7'd113}:		p = 14'd11865;
            {7'd105,7'd114}:		p = 14'd11970;
            {7'd105,7'd115}:		p = 14'd12075;
            {7'd105,7'd116}:		p = 14'd12180;
            {7'd105,7'd117}:		p = 14'd12285;
            {7'd105,7'd118}:		p = 14'd12390;
            {7'd105,7'd119}:		p = 14'd12495;
            {7'd105,7'd120}:		p = 14'd12600;
            {7'd105,7'd121}:		p = 14'd12705;
            {7'd105,7'd122}:		p = 14'd12810;
            {7'd105,7'd123}:		p = 14'd12915;
            {7'd105,7'd124}:		p = 14'd13020;
            {7'd105,7'd125}:		p = 14'd13125;
            {7'd105,7'd126}:		p = 14'd13230;
            {7'd105,7'd127}:		p = 14'd13335;
            {7'd106,7'd0}:		p = 14'd0;
            {7'd106,7'd1}:		p = 14'd106;
            {7'd106,7'd2}:		p = 14'd212;
            {7'd106,7'd3}:		p = 14'd318;
            {7'd106,7'd4}:		p = 14'd424;
            {7'd106,7'd5}:		p = 14'd530;
            {7'd106,7'd6}:		p = 14'd636;
            {7'd106,7'd7}:		p = 14'd742;
            {7'd106,7'd8}:		p = 14'd848;
            {7'd106,7'd9}:		p = 14'd954;
            {7'd106,7'd10}:		p = 14'd1060;
            {7'd106,7'd11}:		p = 14'd1166;
            {7'd106,7'd12}:		p = 14'd1272;
            {7'd106,7'd13}:		p = 14'd1378;
            {7'd106,7'd14}:		p = 14'd1484;
            {7'd106,7'd15}:		p = 14'd1590;
            {7'd106,7'd16}:		p = 14'd1696;
            {7'd106,7'd17}:		p = 14'd1802;
            {7'd106,7'd18}:		p = 14'd1908;
            {7'd106,7'd19}:		p = 14'd2014;
            {7'd106,7'd20}:		p = 14'd2120;
            {7'd106,7'd21}:		p = 14'd2226;
            {7'd106,7'd22}:		p = 14'd2332;
            {7'd106,7'd23}:		p = 14'd2438;
            {7'd106,7'd24}:		p = 14'd2544;
            {7'd106,7'd25}:		p = 14'd2650;
            {7'd106,7'd26}:		p = 14'd2756;
            {7'd106,7'd27}:		p = 14'd2862;
            {7'd106,7'd28}:		p = 14'd2968;
            {7'd106,7'd29}:		p = 14'd3074;
            {7'd106,7'd30}:		p = 14'd3180;
            {7'd106,7'd31}:		p = 14'd3286;
            {7'd106,7'd32}:		p = 14'd3392;
            {7'd106,7'd33}:		p = 14'd3498;
            {7'd106,7'd34}:		p = 14'd3604;
            {7'd106,7'd35}:		p = 14'd3710;
            {7'd106,7'd36}:		p = 14'd3816;
            {7'd106,7'd37}:		p = 14'd3922;
            {7'd106,7'd38}:		p = 14'd4028;
            {7'd106,7'd39}:		p = 14'd4134;
            {7'd106,7'd40}:		p = 14'd4240;
            {7'd106,7'd41}:		p = 14'd4346;
            {7'd106,7'd42}:		p = 14'd4452;
            {7'd106,7'd43}:		p = 14'd4558;
            {7'd106,7'd44}:		p = 14'd4664;
            {7'd106,7'd45}:		p = 14'd4770;
            {7'd106,7'd46}:		p = 14'd4876;
            {7'd106,7'd47}:		p = 14'd4982;
            {7'd106,7'd48}:		p = 14'd5088;
            {7'd106,7'd49}:		p = 14'd5194;
            {7'd106,7'd50}:		p = 14'd5300;
            {7'd106,7'd51}:		p = 14'd5406;
            {7'd106,7'd52}:		p = 14'd5512;
            {7'd106,7'd53}:		p = 14'd5618;
            {7'd106,7'd54}:		p = 14'd5724;
            {7'd106,7'd55}:		p = 14'd5830;
            {7'd106,7'd56}:		p = 14'd5936;
            {7'd106,7'd57}:		p = 14'd6042;
            {7'd106,7'd58}:		p = 14'd6148;
            {7'd106,7'd59}:		p = 14'd6254;
            {7'd106,7'd60}:		p = 14'd6360;
            {7'd106,7'd61}:		p = 14'd6466;
            {7'd106,7'd62}:		p = 14'd6572;
            {7'd106,7'd63}:		p = 14'd6678;
            {7'd106,7'd64}:		p = 14'd6784;
            {7'd106,7'd65}:		p = 14'd6890;
            {7'd106,7'd66}:		p = 14'd6996;
            {7'd106,7'd67}:		p = 14'd7102;
            {7'd106,7'd68}:		p = 14'd7208;
            {7'd106,7'd69}:		p = 14'd7314;
            {7'd106,7'd70}:		p = 14'd7420;
            {7'd106,7'd71}:		p = 14'd7526;
            {7'd106,7'd72}:		p = 14'd7632;
            {7'd106,7'd73}:		p = 14'd7738;
            {7'd106,7'd74}:		p = 14'd7844;
            {7'd106,7'd75}:		p = 14'd7950;
            {7'd106,7'd76}:		p = 14'd8056;
            {7'd106,7'd77}:		p = 14'd8162;
            {7'd106,7'd78}:		p = 14'd8268;
            {7'd106,7'd79}:		p = 14'd8374;
            {7'd106,7'd80}:		p = 14'd8480;
            {7'd106,7'd81}:		p = 14'd8586;
            {7'd106,7'd82}:		p = 14'd8692;
            {7'd106,7'd83}:		p = 14'd8798;
            {7'd106,7'd84}:		p = 14'd8904;
            {7'd106,7'd85}:		p = 14'd9010;
            {7'd106,7'd86}:		p = 14'd9116;
            {7'd106,7'd87}:		p = 14'd9222;
            {7'd106,7'd88}:		p = 14'd9328;
            {7'd106,7'd89}:		p = 14'd9434;
            {7'd106,7'd90}:		p = 14'd9540;
            {7'd106,7'd91}:		p = 14'd9646;
            {7'd106,7'd92}:		p = 14'd9752;
            {7'd106,7'd93}:		p = 14'd9858;
            {7'd106,7'd94}:		p = 14'd9964;
            {7'd106,7'd95}:		p = 14'd10070;
            {7'd106,7'd96}:		p = 14'd10176;
            {7'd106,7'd97}:		p = 14'd10282;
            {7'd106,7'd98}:		p = 14'd10388;
            {7'd106,7'd99}:		p = 14'd10494;
            {7'd106,7'd100}:		p = 14'd10600;
            {7'd106,7'd101}:		p = 14'd10706;
            {7'd106,7'd102}:		p = 14'd10812;
            {7'd106,7'd103}:		p = 14'd10918;
            {7'd106,7'd104}:		p = 14'd11024;
            {7'd106,7'd105}:		p = 14'd11130;
            {7'd106,7'd106}:		p = 14'd11236;
            {7'd106,7'd107}:		p = 14'd11342;
            {7'd106,7'd108}:		p = 14'd11448;
            {7'd106,7'd109}:		p = 14'd11554;
            {7'd106,7'd110}:		p = 14'd11660;
            {7'd106,7'd111}:		p = 14'd11766;
            {7'd106,7'd112}:		p = 14'd11872;
            {7'd106,7'd113}:		p = 14'd11978;
            {7'd106,7'd114}:		p = 14'd12084;
            {7'd106,7'd115}:		p = 14'd12190;
            {7'd106,7'd116}:		p = 14'd12296;
            {7'd106,7'd117}:		p = 14'd12402;
            {7'd106,7'd118}:		p = 14'd12508;
            {7'd106,7'd119}:		p = 14'd12614;
            {7'd106,7'd120}:		p = 14'd12720;
            {7'd106,7'd121}:		p = 14'd12826;
            {7'd106,7'd122}:		p = 14'd12932;
            {7'd106,7'd123}:		p = 14'd13038;
            {7'd106,7'd124}:		p = 14'd13144;
            {7'd106,7'd125}:		p = 14'd13250;
            {7'd106,7'd126}:		p = 14'd13356;
            {7'd106,7'd127}:		p = 14'd13462;
            {7'd107,7'd0}:		p = 14'd0;
            {7'd107,7'd1}:		p = 14'd107;
            {7'd107,7'd2}:		p = 14'd214;
            {7'd107,7'd3}:		p = 14'd321;
            {7'd107,7'd4}:		p = 14'd428;
            {7'd107,7'd5}:		p = 14'd535;
            {7'd107,7'd6}:		p = 14'd642;
            {7'd107,7'd7}:		p = 14'd749;
            {7'd107,7'd8}:		p = 14'd856;
            {7'd107,7'd9}:		p = 14'd963;
            {7'd107,7'd10}:		p = 14'd1070;
            {7'd107,7'd11}:		p = 14'd1177;
            {7'd107,7'd12}:		p = 14'd1284;
            {7'd107,7'd13}:		p = 14'd1391;
            {7'd107,7'd14}:		p = 14'd1498;
            {7'd107,7'd15}:		p = 14'd1605;
            {7'd107,7'd16}:		p = 14'd1712;
            {7'd107,7'd17}:		p = 14'd1819;
            {7'd107,7'd18}:		p = 14'd1926;
            {7'd107,7'd19}:		p = 14'd2033;
            {7'd107,7'd20}:		p = 14'd2140;
            {7'd107,7'd21}:		p = 14'd2247;
            {7'd107,7'd22}:		p = 14'd2354;
            {7'd107,7'd23}:		p = 14'd2461;
            {7'd107,7'd24}:		p = 14'd2568;
            {7'd107,7'd25}:		p = 14'd2675;
            {7'd107,7'd26}:		p = 14'd2782;
            {7'd107,7'd27}:		p = 14'd2889;
            {7'd107,7'd28}:		p = 14'd2996;
            {7'd107,7'd29}:		p = 14'd3103;
            {7'd107,7'd30}:		p = 14'd3210;
            {7'd107,7'd31}:		p = 14'd3317;
            {7'd107,7'd32}:		p = 14'd3424;
            {7'd107,7'd33}:		p = 14'd3531;
            {7'd107,7'd34}:		p = 14'd3638;
            {7'd107,7'd35}:		p = 14'd3745;
            {7'd107,7'd36}:		p = 14'd3852;
            {7'd107,7'd37}:		p = 14'd3959;
            {7'd107,7'd38}:		p = 14'd4066;
            {7'd107,7'd39}:		p = 14'd4173;
            {7'd107,7'd40}:		p = 14'd4280;
            {7'd107,7'd41}:		p = 14'd4387;
            {7'd107,7'd42}:		p = 14'd4494;
            {7'd107,7'd43}:		p = 14'd4601;
            {7'd107,7'd44}:		p = 14'd4708;
            {7'd107,7'd45}:		p = 14'd4815;
            {7'd107,7'd46}:		p = 14'd4922;
            {7'd107,7'd47}:		p = 14'd5029;
            {7'd107,7'd48}:		p = 14'd5136;
            {7'd107,7'd49}:		p = 14'd5243;
            {7'd107,7'd50}:		p = 14'd5350;
            {7'd107,7'd51}:		p = 14'd5457;
            {7'd107,7'd52}:		p = 14'd5564;
            {7'd107,7'd53}:		p = 14'd5671;
            {7'd107,7'd54}:		p = 14'd5778;
            {7'd107,7'd55}:		p = 14'd5885;
            {7'd107,7'd56}:		p = 14'd5992;
            {7'd107,7'd57}:		p = 14'd6099;
            {7'd107,7'd58}:		p = 14'd6206;
            {7'd107,7'd59}:		p = 14'd6313;
            {7'd107,7'd60}:		p = 14'd6420;
            {7'd107,7'd61}:		p = 14'd6527;
            {7'd107,7'd62}:		p = 14'd6634;
            {7'd107,7'd63}:		p = 14'd6741;
            {7'd107,7'd64}:		p = 14'd6848;
            {7'd107,7'd65}:		p = 14'd6955;
            {7'd107,7'd66}:		p = 14'd7062;
            {7'd107,7'd67}:		p = 14'd7169;
            {7'd107,7'd68}:		p = 14'd7276;
            {7'd107,7'd69}:		p = 14'd7383;
            {7'd107,7'd70}:		p = 14'd7490;
            {7'd107,7'd71}:		p = 14'd7597;
            {7'd107,7'd72}:		p = 14'd7704;
            {7'd107,7'd73}:		p = 14'd7811;
            {7'd107,7'd74}:		p = 14'd7918;
            {7'd107,7'd75}:		p = 14'd8025;
            {7'd107,7'd76}:		p = 14'd8132;
            {7'd107,7'd77}:		p = 14'd8239;
            {7'd107,7'd78}:		p = 14'd8346;
            {7'd107,7'd79}:		p = 14'd8453;
            {7'd107,7'd80}:		p = 14'd8560;
            {7'd107,7'd81}:		p = 14'd8667;
            {7'd107,7'd82}:		p = 14'd8774;
            {7'd107,7'd83}:		p = 14'd8881;
            {7'd107,7'd84}:		p = 14'd8988;
            {7'd107,7'd85}:		p = 14'd9095;
            {7'd107,7'd86}:		p = 14'd9202;
            {7'd107,7'd87}:		p = 14'd9309;
            {7'd107,7'd88}:		p = 14'd9416;
            {7'd107,7'd89}:		p = 14'd9523;
            {7'd107,7'd90}:		p = 14'd9630;
            {7'd107,7'd91}:		p = 14'd9737;
            {7'd107,7'd92}:		p = 14'd9844;
            {7'd107,7'd93}:		p = 14'd9951;
            {7'd107,7'd94}:		p = 14'd10058;
            {7'd107,7'd95}:		p = 14'd10165;
            {7'd107,7'd96}:		p = 14'd10272;
            {7'd107,7'd97}:		p = 14'd10379;
            {7'd107,7'd98}:		p = 14'd10486;
            {7'd107,7'd99}:		p = 14'd10593;
            {7'd107,7'd100}:		p = 14'd10700;
            {7'd107,7'd101}:		p = 14'd10807;
            {7'd107,7'd102}:		p = 14'd10914;
            {7'd107,7'd103}:		p = 14'd11021;
            {7'd107,7'd104}:		p = 14'd11128;
            {7'd107,7'd105}:		p = 14'd11235;
            {7'd107,7'd106}:		p = 14'd11342;
            {7'd107,7'd107}:		p = 14'd11449;
            {7'd107,7'd108}:		p = 14'd11556;
            {7'd107,7'd109}:		p = 14'd11663;
            {7'd107,7'd110}:		p = 14'd11770;
            {7'd107,7'd111}:		p = 14'd11877;
            {7'd107,7'd112}:		p = 14'd11984;
            {7'd107,7'd113}:		p = 14'd12091;
            {7'd107,7'd114}:		p = 14'd12198;
            {7'd107,7'd115}:		p = 14'd12305;
            {7'd107,7'd116}:		p = 14'd12412;
            {7'd107,7'd117}:		p = 14'd12519;
            {7'd107,7'd118}:		p = 14'd12626;
            {7'd107,7'd119}:		p = 14'd12733;
            {7'd107,7'd120}:		p = 14'd12840;
            {7'd107,7'd121}:		p = 14'd12947;
            {7'd107,7'd122}:		p = 14'd13054;
            {7'd107,7'd123}:		p = 14'd13161;
            {7'd107,7'd124}:		p = 14'd13268;
            {7'd107,7'd125}:		p = 14'd13375;
            {7'd107,7'd126}:		p = 14'd13482;
            {7'd107,7'd127}:		p = 14'd13589;
            {7'd108,7'd0}:		p = 14'd0;
            {7'd108,7'd1}:		p = 14'd108;
            {7'd108,7'd2}:		p = 14'd216;
            {7'd108,7'd3}:		p = 14'd324;
            {7'd108,7'd4}:		p = 14'd432;
            {7'd108,7'd5}:		p = 14'd540;
            {7'd108,7'd6}:		p = 14'd648;
            {7'd108,7'd7}:		p = 14'd756;
            {7'd108,7'd8}:		p = 14'd864;
            {7'd108,7'd9}:		p = 14'd972;
            {7'd108,7'd10}:		p = 14'd1080;
            {7'd108,7'd11}:		p = 14'd1188;
            {7'd108,7'd12}:		p = 14'd1296;
            {7'd108,7'd13}:		p = 14'd1404;
            {7'd108,7'd14}:		p = 14'd1512;
            {7'd108,7'd15}:		p = 14'd1620;
            {7'd108,7'd16}:		p = 14'd1728;
            {7'd108,7'd17}:		p = 14'd1836;
            {7'd108,7'd18}:		p = 14'd1944;
            {7'd108,7'd19}:		p = 14'd2052;
            {7'd108,7'd20}:		p = 14'd2160;
            {7'd108,7'd21}:		p = 14'd2268;
            {7'd108,7'd22}:		p = 14'd2376;
            {7'd108,7'd23}:		p = 14'd2484;
            {7'd108,7'd24}:		p = 14'd2592;
            {7'd108,7'd25}:		p = 14'd2700;
            {7'd108,7'd26}:		p = 14'd2808;
            {7'd108,7'd27}:		p = 14'd2916;
            {7'd108,7'd28}:		p = 14'd3024;
            {7'd108,7'd29}:		p = 14'd3132;
            {7'd108,7'd30}:		p = 14'd3240;
            {7'd108,7'd31}:		p = 14'd3348;
            {7'd108,7'd32}:		p = 14'd3456;
            {7'd108,7'd33}:		p = 14'd3564;
            {7'd108,7'd34}:		p = 14'd3672;
            {7'd108,7'd35}:		p = 14'd3780;
            {7'd108,7'd36}:		p = 14'd3888;
            {7'd108,7'd37}:		p = 14'd3996;
            {7'd108,7'd38}:		p = 14'd4104;
            {7'd108,7'd39}:		p = 14'd4212;
            {7'd108,7'd40}:		p = 14'd4320;
            {7'd108,7'd41}:		p = 14'd4428;
            {7'd108,7'd42}:		p = 14'd4536;
            {7'd108,7'd43}:		p = 14'd4644;
            {7'd108,7'd44}:		p = 14'd4752;
            {7'd108,7'd45}:		p = 14'd4860;
            {7'd108,7'd46}:		p = 14'd4968;
            {7'd108,7'd47}:		p = 14'd5076;
            {7'd108,7'd48}:		p = 14'd5184;
            {7'd108,7'd49}:		p = 14'd5292;
            {7'd108,7'd50}:		p = 14'd5400;
            {7'd108,7'd51}:		p = 14'd5508;
            {7'd108,7'd52}:		p = 14'd5616;
            {7'd108,7'd53}:		p = 14'd5724;
            {7'd108,7'd54}:		p = 14'd5832;
            {7'd108,7'd55}:		p = 14'd5940;
            {7'd108,7'd56}:		p = 14'd6048;
            {7'd108,7'd57}:		p = 14'd6156;
            {7'd108,7'd58}:		p = 14'd6264;
            {7'd108,7'd59}:		p = 14'd6372;
            {7'd108,7'd60}:		p = 14'd6480;
            {7'd108,7'd61}:		p = 14'd6588;
            {7'd108,7'd62}:		p = 14'd6696;
            {7'd108,7'd63}:		p = 14'd6804;
            {7'd108,7'd64}:		p = 14'd6912;
            {7'd108,7'd65}:		p = 14'd7020;
            {7'd108,7'd66}:		p = 14'd7128;
            {7'd108,7'd67}:		p = 14'd7236;
            {7'd108,7'd68}:		p = 14'd7344;
            {7'd108,7'd69}:		p = 14'd7452;
            {7'd108,7'd70}:		p = 14'd7560;
            {7'd108,7'd71}:		p = 14'd7668;
            {7'd108,7'd72}:		p = 14'd7776;
            {7'd108,7'd73}:		p = 14'd7884;
            {7'd108,7'd74}:		p = 14'd7992;
            {7'd108,7'd75}:		p = 14'd8100;
            {7'd108,7'd76}:		p = 14'd8208;
            {7'd108,7'd77}:		p = 14'd8316;
            {7'd108,7'd78}:		p = 14'd8424;
            {7'd108,7'd79}:		p = 14'd8532;
            {7'd108,7'd80}:		p = 14'd8640;
            {7'd108,7'd81}:		p = 14'd8748;
            {7'd108,7'd82}:		p = 14'd8856;
            {7'd108,7'd83}:		p = 14'd8964;
            {7'd108,7'd84}:		p = 14'd9072;
            {7'd108,7'd85}:		p = 14'd9180;
            {7'd108,7'd86}:		p = 14'd9288;
            {7'd108,7'd87}:		p = 14'd9396;
            {7'd108,7'd88}:		p = 14'd9504;
            {7'd108,7'd89}:		p = 14'd9612;
            {7'd108,7'd90}:		p = 14'd9720;
            {7'd108,7'd91}:		p = 14'd9828;
            {7'd108,7'd92}:		p = 14'd9936;
            {7'd108,7'd93}:		p = 14'd10044;
            {7'd108,7'd94}:		p = 14'd10152;
            {7'd108,7'd95}:		p = 14'd10260;
            {7'd108,7'd96}:		p = 14'd10368;
            {7'd108,7'd97}:		p = 14'd10476;
            {7'd108,7'd98}:		p = 14'd10584;
            {7'd108,7'd99}:		p = 14'd10692;
            {7'd108,7'd100}:		p = 14'd10800;
            {7'd108,7'd101}:		p = 14'd10908;
            {7'd108,7'd102}:		p = 14'd11016;
            {7'd108,7'd103}:		p = 14'd11124;
            {7'd108,7'd104}:		p = 14'd11232;
            {7'd108,7'd105}:		p = 14'd11340;
            {7'd108,7'd106}:		p = 14'd11448;
            {7'd108,7'd107}:		p = 14'd11556;
            {7'd108,7'd108}:		p = 14'd11664;
            {7'd108,7'd109}:		p = 14'd11772;
            {7'd108,7'd110}:		p = 14'd11880;
            {7'd108,7'd111}:		p = 14'd11988;
            {7'd108,7'd112}:		p = 14'd12096;
            {7'd108,7'd113}:		p = 14'd12204;
            {7'd108,7'd114}:		p = 14'd12312;
            {7'd108,7'd115}:		p = 14'd12420;
            {7'd108,7'd116}:		p = 14'd12528;
            {7'd108,7'd117}:		p = 14'd12636;
            {7'd108,7'd118}:		p = 14'd12744;
            {7'd108,7'd119}:		p = 14'd12852;
            {7'd108,7'd120}:		p = 14'd12960;
            {7'd108,7'd121}:		p = 14'd13068;
            {7'd108,7'd122}:		p = 14'd13176;
            {7'd108,7'd123}:		p = 14'd13284;
            {7'd108,7'd124}:		p = 14'd13392;
            {7'd108,7'd125}:		p = 14'd13500;
            {7'd108,7'd126}:		p = 14'd13608;
            {7'd108,7'd127}:		p = 14'd13716;
            {7'd109,7'd0}:		p = 14'd0;
            {7'd109,7'd1}:		p = 14'd109;
            {7'd109,7'd2}:		p = 14'd218;
            {7'd109,7'd3}:		p = 14'd327;
            {7'd109,7'd4}:		p = 14'd436;
            {7'd109,7'd5}:		p = 14'd545;
            {7'd109,7'd6}:		p = 14'd654;
            {7'd109,7'd7}:		p = 14'd763;
            {7'd109,7'd8}:		p = 14'd872;
            {7'd109,7'd9}:		p = 14'd981;
            {7'd109,7'd10}:		p = 14'd1090;
            {7'd109,7'd11}:		p = 14'd1199;
            {7'd109,7'd12}:		p = 14'd1308;
            {7'd109,7'd13}:		p = 14'd1417;
            {7'd109,7'd14}:		p = 14'd1526;
            {7'd109,7'd15}:		p = 14'd1635;
            {7'd109,7'd16}:		p = 14'd1744;
            {7'd109,7'd17}:		p = 14'd1853;
            {7'd109,7'd18}:		p = 14'd1962;
            {7'd109,7'd19}:		p = 14'd2071;
            {7'd109,7'd20}:		p = 14'd2180;
            {7'd109,7'd21}:		p = 14'd2289;
            {7'd109,7'd22}:		p = 14'd2398;
            {7'd109,7'd23}:		p = 14'd2507;
            {7'd109,7'd24}:		p = 14'd2616;
            {7'd109,7'd25}:		p = 14'd2725;
            {7'd109,7'd26}:		p = 14'd2834;
            {7'd109,7'd27}:		p = 14'd2943;
            {7'd109,7'd28}:		p = 14'd3052;
            {7'd109,7'd29}:		p = 14'd3161;
            {7'd109,7'd30}:		p = 14'd3270;
            {7'd109,7'd31}:		p = 14'd3379;
            {7'd109,7'd32}:		p = 14'd3488;
            {7'd109,7'd33}:		p = 14'd3597;
            {7'd109,7'd34}:		p = 14'd3706;
            {7'd109,7'd35}:		p = 14'd3815;
            {7'd109,7'd36}:		p = 14'd3924;
            {7'd109,7'd37}:		p = 14'd4033;
            {7'd109,7'd38}:		p = 14'd4142;
            {7'd109,7'd39}:		p = 14'd4251;
            {7'd109,7'd40}:		p = 14'd4360;
            {7'd109,7'd41}:		p = 14'd4469;
            {7'd109,7'd42}:		p = 14'd4578;
            {7'd109,7'd43}:		p = 14'd4687;
            {7'd109,7'd44}:		p = 14'd4796;
            {7'd109,7'd45}:		p = 14'd4905;
            {7'd109,7'd46}:		p = 14'd5014;
            {7'd109,7'd47}:		p = 14'd5123;
            {7'd109,7'd48}:		p = 14'd5232;
            {7'd109,7'd49}:		p = 14'd5341;
            {7'd109,7'd50}:		p = 14'd5450;
            {7'd109,7'd51}:		p = 14'd5559;
            {7'd109,7'd52}:		p = 14'd5668;
            {7'd109,7'd53}:		p = 14'd5777;
            {7'd109,7'd54}:		p = 14'd5886;
            {7'd109,7'd55}:		p = 14'd5995;
            {7'd109,7'd56}:		p = 14'd6104;
            {7'd109,7'd57}:		p = 14'd6213;
            {7'd109,7'd58}:		p = 14'd6322;
            {7'd109,7'd59}:		p = 14'd6431;
            {7'd109,7'd60}:		p = 14'd6540;
            {7'd109,7'd61}:		p = 14'd6649;
            {7'd109,7'd62}:		p = 14'd6758;
            {7'd109,7'd63}:		p = 14'd6867;
            {7'd109,7'd64}:		p = 14'd6976;
            {7'd109,7'd65}:		p = 14'd7085;
            {7'd109,7'd66}:		p = 14'd7194;
            {7'd109,7'd67}:		p = 14'd7303;
            {7'd109,7'd68}:		p = 14'd7412;
            {7'd109,7'd69}:		p = 14'd7521;
            {7'd109,7'd70}:		p = 14'd7630;
            {7'd109,7'd71}:		p = 14'd7739;
            {7'd109,7'd72}:		p = 14'd7848;
            {7'd109,7'd73}:		p = 14'd7957;
            {7'd109,7'd74}:		p = 14'd8066;
            {7'd109,7'd75}:		p = 14'd8175;
            {7'd109,7'd76}:		p = 14'd8284;
            {7'd109,7'd77}:		p = 14'd8393;
            {7'd109,7'd78}:		p = 14'd8502;
            {7'd109,7'd79}:		p = 14'd8611;
            {7'd109,7'd80}:		p = 14'd8720;
            {7'd109,7'd81}:		p = 14'd8829;
            {7'd109,7'd82}:		p = 14'd8938;
            {7'd109,7'd83}:		p = 14'd9047;
            {7'd109,7'd84}:		p = 14'd9156;
            {7'd109,7'd85}:		p = 14'd9265;
            {7'd109,7'd86}:		p = 14'd9374;
            {7'd109,7'd87}:		p = 14'd9483;
            {7'd109,7'd88}:		p = 14'd9592;
            {7'd109,7'd89}:		p = 14'd9701;
            {7'd109,7'd90}:		p = 14'd9810;
            {7'd109,7'd91}:		p = 14'd9919;
            {7'd109,7'd92}:		p = 14'd10028;
            {7'd109,7'd93}:		p = 14'd10137;
            {7'd109,7'd94}:		p = 14'd10246;
            {7'd109,7'd95}:		p = 14'd10355;
            {7'd109,7'd96}:		p = 14'd10464;
            {7'd109,7'd97}:		p = 14'd10573;
            {7'd109,7'd98}:		p = 14'd10682;
            {7'd109,7'd99}:		p = 14'd10791;
            {7'd109,7'd100}:		p = 14'd10900;
            {7'd109,7'd101}:		p = 14'd11009;
            {7'd109,7'd102}:		p = 14'd11118;
            {7'd109,7'd103}:		p = 14'd11227;
            {7'd109,7'd104}:		p = 14'd11336;
            {7'd109,7'd105}:		p = 14'd11445;
            {7'd109,7'd106}:		p = 14'd11554;
            {7'd109,7'd107}:		p = 14'd11663;
            {7'd109,7'd108}:		p = 14'd11772;
            {7'd109,7'd109}:		p = 14'd11881;
            {7'd109,7'd110}:		p = 14'd11990;
            {7'd109,7'd111}:		p = 14'd12099;
            {7'd109,7'd112}:		p = 14'd12208;
            {7'd109,7'd113}:		p = 14'd12317;
            {7'd109,7'd114}:		p = 14'd12426;
            {7'd109,7'd115}:		p = 14'd12535;
            {7'd109,7'd116}:		p = 14'd12644;
            {7'd109,7'd117}:		p = 14'd12753;
            {7'd109,7'd118}:		p = 14'd12862;
            {7'd109,7'd119}:		p = 14'd12971;
            {7'd109,7'd120}:		p = 14'd13080;
            {7'd109,7'd121}:		p = 14'd13189;
            {7'd109,7'd122}:		p = 14'd13298;
            {7'd109,7'd123}:		p = 14'd13407;
            {7'd109,7'd124}:		p = 14'd13516;
            {7'd109,7'd125}:		p = 14'd13625;
            {7'd109,7'd126}:		p = 14'd13734;
            {7'd109,7'd127}:		p = 14'd13843;
            {7'd110,7'd0}:		p = 14'd0;
            {7'd110,7'd1}:		p = 14'd110;
            {7'd110,7'd2}:		p = 14'd220;
            {7'd110,7'd3}:		p = 14'd330;
            {7'd110,7'd4}:		p = 14'd440;
            {7'd110,7'd5}:		p = 14'd550;
            {7'd110,7'd6}:		p = 14'd660;
            {7'd110,7'd7}:		p = 14'd770;
            {7'd110,7'd8}:		p = 14'd880;
            {7'd110,7'd9}:		p = 14'd990;
            {7'd110,7'd10}:		p = 14'd1100;
            {7'd110,7'd11}:		p = 14'd1210;
            {7'd110,7'd12}:		p = 14'd1320;
            {7'd110,7'd13}:		p = 14'd1430;
            {7'd110,7'd14}:		p = 14'd1540;
            {7'd110,7'd15}:		p = 14'd1650;
            {7'd110,7'd16}:		p = 14'd1760;
            {7'd110,7'd17}:		p = 14'd1870;
            {7'd110,7'd18}:		p = 14'd1980;
            {7'd110,7'd19}:		p = 14'd2090;
            {7'd110,7'd20}:		p = 14'd2200;
            {7'd110,7'd21}:		p = 14'd2310;
            {7'd110,7'd22}:		p = 14'd2420;
            {7'd110,7'd23}:		p = 14'd2530;
            {7'd110,7'd24}:		p = 14'd2640;
            {7'd110,7'd25}:		p = 14'd2750;
            {7'd110,7'd26}:		p = 14'd2860;
            {7'd110,7'd27}:		p = 14'd2970;
            {7'd110,7'd28}:		p = 14'd3080;
            {7'd110,7'd29}:		p = 14'd3190;
            {7'd110,7'd30}:		p = 14'd3300;
            {7'd110,7'd31}:		p = 14'd3410;
            {7'd110,7'd32}:		p = 14'd3520;
            {7'd110,7'd33}:		p = 14'd3630;
            {7'd110,7'd34}:		p = 14'd3740;
            {7'd110,7'd35}:		p = 14'd3850;
            {7'd110,7'd36}:		p = 14'd3960;
            {7'd110,7'd37}:		p = 14'd4070;
            {7'd110,7'd38}:		p = 14'd4180;
            {7'd110,7'd39}:		p = 14'd4290;
            {7'd110,7'd40}:		p = 14'd4400;
            {7'd110,7'd41}:		p = 14'd4510;
            {7'd110,7'd42}:		p = 14'd4620;
            {7'd110,7'd43}:		p = 14'd4730;
            {7'd110,7'd44}:		p = 14'd4840;
            {7'd110,7'd45}:		p = 14'd4950;
            {7'd110,7'd46}:		p = 14'd5060;
            {7'd110,7'd47}:		p = 14'd5170;
            {7'd110,7'd48}:		p = 14'd5280;
            {7'd110,7'd49}:		p = 14'd5390;
            {7'd110,7'd50}:		p = 14'd5500;
            {7'd110,7'd51}:		p = 14'd5610;
            {7'd110,7'd52}:		p = 14'd5720;
            {7'd110,7'd53}:		p = 14'd5830;
            {7'd110,7'd54}:		p = 14'd5940;
            {7'd110,7'd55}:		p = 14'd6050;
            {7'd110,7'd56}:		p = 14'd6160;
            {7'd110,7'd57}:		p = 14'd6270;
            {7'd110,7'd58}:		p = 14'd6380;
            {7'd110,7'd59}:		p = 14'd6490;
            {7'd110,7'd60}:		p = 14'd6600;
            {7'd110,7'd61}:		p = 14'd6710;
            {7'd110,7'd62}:		p = 14'd6820;
            {7'd110,7'd63}:		p = 14'd6930;
            {7'd110,7'd64}:		p = 14'd7040;
            {7'd110,7'd65}:		p = 14'd7150;
            {7'd110,7'd66}:		p = 14'd7260;
            {7'd110,7'd67}:		p = 14'd7370;
            {7'd110,7'd68}:		p = 14'd7480;
            {7'd110,7'd69}:		p = 14'd7590;
            {7'd110,7'd70}:		p = 14'd7700;
            {7'd110,7'd71}:		p = 14'd7810;
            {7'd110,7'd72}:		p = 14'd7920;
            {7'd110,7'd73}:		p = 14'd8030;
            {7'd110,7'd74}:		p = 14'd8140;
            {7'd110,7'd75}:		p = 14'd8250;
            {7'd110,7'd76}:		p = 14'd8360;
            {7'd110,7'd77}:		p = 14'd8470;
            {7'd110,7'd78}:		p = 14'd8580;
            {7'd110,7'd79}:		p = 14'd8690;
            {7'd110,7'd80}:		p = 14'd8800;
            {7'd110,7'd81}:		p = 14'd8910;
            {7'd110,7'd82}:		p = 14'd9020;
            {7'd110,7'd83}:		p = 14'd9130;
            {7'd110,7'd84}:		p = 14'd9240;
            {7'd110,7'd85}:		p = 14'd9350;
            {7'd110,7'd86}:		p = 14'd9460;
            {7'd110,7'd87}:		p = 14'd9570;
            {7'd110,7'd88}:		p = 14'd9680;
            {7'd110,7'd89}:		p = 14'd9790;
            {7'd110,7'd90}:		p = 14'd9900;
            {7'd110,7'd91}:		p = 14'd10010;
            {7'd110,7'd92}:		p = 14'd10120;
            {7'd110,7'd93}:		p = 14'd10230;
            {7'd110,7'd94}:		p = 14'd10340;
            {7'd110,7'd95}:		p = 14'd10450;
            {7'd110,7'd96}:		p = 14'd10560;
            {7'd110,7'd97}:		p = 14'd10670;
            {7'd110,7'd98}:		p = 14'd10780;
            {7'd110,7'd99}:		p = 14'd10890;
            {7'd110,7'd100}:		p = 14'd11000;
            {7'd110,7'd101}:		p = 14'd11110;
            {7'd110,7'd102}:		p = 14'd11220;
            {7'd110,7'd103}:		p = 14'd11330;
            {7'd110,7'd104}:		p = 14'd11440;
            {7'd110,7'd105}:		p = 14'd11550;
            {7'd110,7'd106}:		p = 14'd11660;
            {7'd110,7'd107}:		p = 14'd11770;
            {7'd110,7'd108}:		p = 14'd11880;
            {7'd110,7'd109}:		p = 14'd11990;
            {7'd110,7'd110}:		p = 14'd12100;
            {7'd110,7'd111}:		p = 14'd12210;
            {7'd110,7'd112}:		p = 14'd12320;
            {7'd110,7'd113}:		p = 14'd12430;
            {7'd110,7'd114}:		p = 14'd12540;
            {7'd110,7'd115}:		p = 14'd12650;
            {7'd110,7'd116}:		p = 14'd12760;
            {7'd110,7'd117}:		p = 14'd12870;
            {7'd110,7'd118}:		p = 14'd12980;
            {7'd110,7'd119}:		p = 14'd13090;
            {7'd110,7'd120}:		p = 14'd13200;
            {7'd110,7'd121}:		p = 14'd13310;
            {7'd110,7'd122}:		p = 14'd13420;
            {7'd110,7'd123}:		p = 14'd13530;
            {7'd110,7'd124}:		p = 14'd13640;
            {7'd110,7'd125}:		p = 14'd13750;
            {7'd110,7'd126}:		p = 14'd13860;
            {7'd110,7'd127}:		p = 14'd13970;
            {7'd111,7'd0}:		p = 14'd0;
            {7'd111,7'd1}:		p = 14'd111;
            {7'd111,7'd2}:		p = 14'd222;
            {7'd111,7'd3}:		p = 14'd333;
            {7'd111,7'd4}:		p = 14'd444;
            {7'd111,7'd5}:		p = 14'd555;
            {7'd111,7'd6}:		p = 14'd666;
            {7'd111,7'd7}:		p = 14'd777;
            {7'd111,7'd8}:		p = 14'd888;
            {7'd111,7'd9}:		p = 14'd999;
            {7'd111,7'd10}:		p = 14'd1110;
            {7'd111,7'd11}:		p = 14'd1221;
            {7'd111,7'd12}:		p = 14'd1332;
            {7'd111,7'd13}:		p = 14'd1443;
            {7'd111,7'd14}:		p = 14'd1554;
            {7'd111,7'd15}:		p = 14'd1665;
            {7'd111,7'd16}:		p = 14'd1776;
            {7'd111,7'd17}:		p = 14'd1887;
            {7'd111,7'd18}:		p = 14'd1998;
            {7'd111,7'd19}:		p = 14'd2109;
            {7'd111,7'd20}:		p = 14'd2220;
            {7'd111,7'd21}:		p = 14'd2331;
            {7'd111,7'd22}:		p = 14'd2442;
            {7'd111,7'd23}:		p = 14'd2553;
            {7'd111,7'd24}:		p = 14'd2664;
            {7'd111,7'd25}:		p = 14'd2775;
            {7'd111,7'd26}:		p = 14'd2886;
            {7'd111,7'd27}:		p = 14'd2997;
            {7'd111,7'd28}:		p = 14'd3108;
            {7'd111,7'd29}:		p = 14'd3219;
            {7'd111,7'd30}:		p = 14'd3330;
            {7'd111,7'd31}:		p = 14'd3441;
            {7'd111,7'd32}:		p = 14'd3552;
            {7'd111,7'd33}:		p = 14'd3663;
            {7'd111,7'd34}:		p = 14'd3774;
            {7'd111,7'd35}:		p = 14'd3885;
            {7'd111,7'd36}:		p = 14'd3996;
            {7'd111,7'd37}:		p = 14'd4107;
            {7'd111,7'd38}:		p = 14'd4218;
            {7'd111,7'd39}:		p = 14'd4329;
            {7'd111,7'd40}:		p = 14'd4440;
            {7'd111,7'd41}:		p = 14'd4551;
            {7'd111,7'd42}:		p = 14'd4662;
            {7'd111,7'd43}:		p = 14'd4773;
            {7'd111,7'd44}:		p = 14'd4884;
            {7'd111,7'd45}:		p = 14'd4995;
            {7'd111,7'd46}:		p = 14'd5106;
            {7'd111,7'd47}:		p = 14'd5217;
            {7'd111,7'd48}:		p = 14'd5328;
            {7'd111,7'd49}:		p = 14'd5439;
            {7'd111,7'd50}:		p = 14'd5550;
            {7'd111,7'd51}:		p = 14'd5661;
            {7'd111,7'd52}:		p = 14'd5772;
            {7'd111,7'd53}:		p = 14'd5883;
            {7'd111,7'd54}:		p = 14'd5994;
            {7'd111,7'd55}:		p = 14'd6105;
            {7'd111,7'd56}:		p = 14'd6216;
            {7'd111,7'd57}:		p = 14'd6327;
            {7'd111,7'd58}:		p = 14'd6438;
            {7'd111,7'd59}:		p = 14'd6549;
            {7'd111,7'd60}:		p = 14'd6660;
            {7'd111,7'd61}:		p = 14'd6771;
            {7'd111,7'd62}:		p = 14'd6882;
            {7'd111,7'd63}:		p = 14'd6993;
            {7'd111,7'd64}:		p = 14'd7104;
            {7'd111,7'd65}:		p = 14'd7215;
            {7'd111,7'd66}:		p = 14'd7326;
            {7'd111,7'd67}:		p = 14'd7437;
            {7'd111,7'd68}:		p = 14'd7548;
            {7'd111,7'd69}:		p = 14'd7659;
            {7'd111,7'd70}:		p = 14'd7770;
            {7'd111,7'd71}:		p = 14'd7881;
            {7'd111,7'd72}:		p = 14'd7992;
            {7'd111,7'd73}:		p = 14'd8103;
            {7'd111,7'd74}:		p = 14'd8214;
            {7'd111,7'd75}:		p = 14'd8325;
            {7'd111,7'd76}:		p = 14'd8436;
            {7'd111,7'd77}:		p = 14'd8547;
            {7'd111,7'd78}:		p = 14'd8658;
            {7'd111,7'd79}:		p = 14'd8769;
            {7'd111,7'd80}:		p = 14'd8880;
            {7'd111,7'd81}:		p = 14'd8991;
            {7'd111,7'd82}:		p = 14'd9102;
            {7'd111,7'd83}:		p = 14'd9213;
            {7'd111,7'd84}:		p = 14'd9324;
            {7'd111,7'd85}:		p = 14'd9435;
            {7'd111,7'd86}:		p = 14'd9546;
            {7'd111,7'd87}:		p = 14'd9657;
            {7'd111,7'd88}:		p = 14'd9768;
            {7'd111,7'd89}:		p = 14'd9879;
            {7'd111,7'd90}:		p = 14'd9990;
            {7'd111,7'd91}:		p = 14'd10101;
            {7'd111,7'd92}:		p = 14'd10212;
            {7'd111,7'd93}:		p = 14'd10323;
            {7'd111,7'd94}:		p = 14'd10434;
            {7'd111,7'd95}:		p = 14'd10545;
            {7'd111,7'd96}:		p = 14'd10656;
            {7'd111,7'd97}:		p = 14'd10767;
            {7'd111,7'd98}:		p = 14'd10878;
            {7'd111,7'd99}:		p = 14'd10989;
            {7'd111,7'd100}:		p = 14'd11100;
            {7'd111,7'd101}:		p = 14'd11211;
            {7'd111,7'd102}:		p = 14'd11322;
            {7'd111,7'd103}:		p = 14'd11433;
            {7'd111,7'd104}:		p = 14'd11544;
            {7'd111,7'd105}:		p = 14'd11655;
            {7'd111,7'd106}:		p = 14'd11766;
            {7'd111,7'd107}:		p = 14'd11877;
            {7'd111,7'd108}:		p = 14'd11988;
            {7'd111,7'd109}:		p = 14'd12099;
            {7'd111,7'd110}:		p = 14'd12210;
            {7'd111,7'd111}:		p = 14'd12321;
            {7'd111,7'd112}:		p = 14'd12432;
            {7'd111,7'd113}:		p = 14'd12543;
            {7'd111,7'd114}:		p = 14'd12654;
            {7'd111,7'd115}:		p = 14'd12765;
            {7'd111,7'd116}:		p = 14'd12876;
            {7'd111,7'd117}:		p = 14'd12987;
            {7'd111,7'd118}:		p = 14'd13098;
            {7'd111,7'd119}:		p = 14'd13209;
            {7'd111,7'd120}:		p = 14'd13320;
            {7'd111,7'd121}:		p = 14'd13431;
            {7'd111,7'd122}:		p = 14'd13542;
            {7'd111,7'd123}:		p = 14'd13653;
            {7'd111,7'd124}:		p = 14'd13764;
            {7'd111,7'd125}:		p = 14'd13875;
            {7'd111,7'd126}:		p = 14'd13986;
            {7'd111,7'd127}:		p = 14'd14097;
            {7'd112,7'd0}:		p = 14'd0;
            {7'd112,7'd1}:		p = 14'd112;
            {7'd112,7'd2}:		p = 14'd224;
            {7'd112,7'd3}:		p = 14'd336;
            {7'd112,7'd4}:		p = 14'd448;
            {7'd112,7'd5}:		p = 14'd560;
            {7'd112,7'd6}:		p = 14'd672;
            {7'd112,7'd7}:		p = 14'd784;
            {7'd112,7'd8}:		p = 14'd896;
            {7'd112,7'd9}:		p = 14'd1008;
            {7'd112,7'd10}:		p = 14'd1120;
            {7'd112,7'd11}:		p = 14'd1232;
            {7'd112,7'd12}:		p = 14'd1344;
            {7'd112,7'd13}:		p = 14'd1456;
            {7'd112,7'd14}:		p = 14'd1568;
            {7'd112,7'd15}:		p = 14'd1680;
            {7'd112,7'd16}:		p = 14'd1792;
            {7'd112,7'd17}:		p = 14'd1904;
            {7'd112,7'd18}:		p = 14'd2016;
            {7'd112,7'd19}:		p = 14'd2128;
            {7'd112,7'd20}:		p = 14'd2240;
            {7'd112,7'd21}:		p = 14'd2352;
            {7'd112,7'd22}:		p = 14'd2464;
            {7'd112,7'd23}:		p = 14'd2576;
            {7'd112,7'd24}:		p = 14'd2688;
            {7'd112,7'd25}:		p = 14'd2800;
            {7'd112,7'd26}:		p = 14'd2912;
            {7'd112,7'd27}:		p = 14'd3024;
            {7'd112,7'd28}:		p = 14'd3136;
            {7'd112,7'd29}:		p = 14'd3248;
            {7'd112,7'd30}:		p = 14'd3360;
            {7'd112,7'd31}:		p = 14'd3472;
            {7'd112,7'd32}:		p = 14'd3584;
            {7'd112,7'd33}:		p = 14'd3696;
            {7'd112,7'd34}:		p = 14'd3808;
            {7'd112,7'd35}:		p = 14'd3920;
            {7'd112,7'd36}:		p = 14'd4032;
            {7'd112,7'd37}:		p = 14'd4144;
            {7'd112,7'd38}:		p = 14'd4256;
            {7'd112,7'd39}:		p = 14'd4368;
            {7'd112,7'd40}:		p = 14'd4480;
            {7'd112,7'd41}:		p = 14'd4592;
            {7'd112,7'd42}:		p = 14'd4704;
            {7'd112,7'd43}:		p = 14'd4816;
            {7'd112,7'd44}:		p = 14'd4928;
            {7'd112,7'd45}:		p = 14'd5040;
            {7'd112,7'd46}:		p = 14'd5152;
            {7'd112,7'd47}:		p = 14'd5264;
            {7'd112,7'd48}:		p = 14'd5376;
            {7'd112,7'd49}:		p = 14'd5488;
            {7'd112,7'd50}:		p = 14'd5600;
            {7'd112,7'd51}:		p = 14'd5712;
            {7'd112,7'd52}:		p = 14'd5824;
            {7'd112,7'd53}:		p = 14'd5936;
            {7'd112,7'd54}:		p = 14'd6048;
            {7'd112,7'd55}:		p = 14'd6160;
            {7'd112,7'd56}:		p = 14'd6272;
            {7'd112,7'd57}:		p = 14'd6384;
            {7'd112,7'd58}:		p = 14'd6496;
            {7'd112,7'd59}:		p = 14'd6608;
            {7'd112,7'd60}:		p = 14'd6720;
            {7'd112,7'd61}:		p = 14'd6832;
            {7'd112,7'd62}:		p = 14'd6944;
            {7'd112,7'd63}:		p = 14'd7056;
            {7'd112,7'd64}:		p = 14'd7168;
            {7'd112,7'd65}:		p = 14'd7280;
            {7'd112,7'd66}:		p = 14'd7392;
            {7'd112,7'd67}:		p = 14'd7504;
            {7'd112,7'd68}:		p = 14'd7616;
            {7'd112,7'd69}:		p = 14'd7728;
            {7'd112,7'd70}:		p = 14'd7840;
            {7'd112,7'd71}:		p = 14'd7952;
            {7'd112,7'd72}:		p = 14'd8064;
            {7'd112,7'd73}:		p = 14'd8176;
            {7'd112,7'd74}:		p = 14'd8288;
            {7'd112,7'd75}:		p = 14'd8400;
            {7'd112,7'd76}:		p = 14'd8512;
            {7'd112,7'd77}:		p = 14'd8624;
            {7'd112,7'd78}:		p = 14'd8736;
            {7'd112,7'd79}:		p = 14'd8848;
            {7'd112,7'd80}:		p = 14'd8960;
            {7'd112,7'd81}:		p = 14'd9072;
            {7'd112,7'd82}:		p = 14'd9184;
            {7'd112,7'd83}:		p = 14'd9296;
            {7'd112,7'd84}:		p = 14'd9408;
            {7'd112,7'd85}:		p = 14'd9520;
            {7'd112,7'd86}:		p = 14'd9632;
            {7'd112,7'd87}:		p = 14'd9744;
            {7'd112,7'd88}:		p = 14'd9856;
            {7'd112,7'd89}:		p = 14'd9968;
            {7'd112,7'd90}:		p = 14'd10080;
            {7'd112,7'd91}:		p = 14'd10192;
            {7'd112,7'd92}:		p = 14'd10304;
            {7'd112,7'd93}:		p = 14'd10416;
            {7'd112,7'd94}:		p = 14'd10528;
            {7'd112,7'd95}:		p = 14'd10640;
            {7'd112,7'd96}:		p = 14'd10752;
            {7'd112,7'd97}:		p = 14'd10864;
            {7'd112,7'd98}:		p = 14'd10976;
            {7'd112,7'd99}:		p = 14'd11088;
            {7'd112,7'd100}:		p = 14'd11200;
            {7'd112,7'd101}:		p = 14'd11312;
            {7'd112,7'd102}:		p = 14'd11424;
            {7'd112,7'd103}:		p = 14'd11536;
            {7'd112,7'd104}:		p = 14'd11648;
            {7'd112,7'd105}:		p = 14'd11760;
            {7'd112,7'd106}:		p = 14'd11872;
            {7'd112,7'd107}:		p = 14'd11984;
            {7'd112,7'd108}:		p = 14'd12096;
            {7'd112,7'd109}:		p = 14'd12208;
            {7'd112,7'd110}:		p = 14'd12320;
            {7'd112,7'd111}:		p = 14'd12432;
            {7'd112,7'd112}:		p = 14'd12544;
            {7'd112,7'd113}:		p = 14'd12656;
            {7'd112,7'd114}:		p = 14'd12768;
            {7'd112,7'd115}:		p = 14'd12880;
            {7'd112,7'd116}:		p = 14'd12992;
            {7'd112,7'd117}:		p = 14'd13104;
            {7'd112,7'd118}:		p = 14'd13216;
            {7'd112,7'd119}:		p = 14'd13328;
            {7'd112,7'd120}:		p = 14'd13440;
            {7'd112,7'd121}:		p = 14'd13552;
            {7'd112,7'd122}:		p = 14'd13664;
            {7'd112,7'd123}:		p = 14'd13776;
            {7'd112,7'd124}:		p = 14'd13888;
            {7'd112,7'd125}:		p = 14'd14000;
            {7'd112,7'd126}:		p = 14'd14112;
            {7'd112,7'd127}:		p = 14'd14224;
            {7'd113,7'd0}:		p = 14'd0;
            {7'd113,7'd1}:		p = 14'd113;
            {7'd113,7'd2}:		p = 14'd226;
            {7'd113,7'd3}:		p = 14'd339;
            {7'd113,7'd4}:		p = 14'd452;
            {7'd113,7'd5}:		p = 14'd565;
            {7'd113,7'd6}:		p = 14'd678;
            {7'd113,7'd7}:		p = 14'd791;
            {7'd113,7'd8}:		p = 14'd904;
            {7'd113,7'd9}:		p = 14'd1017;
            {7'd113,7'd10}:		p = 14'd1130;
            {7'd113,7'd11}:		p = 14'd1243;
            {7'd113,7'd12}:		p = 14'd1356;
            {7'd113,7'd13}:		p = 14'd1469;
            {7'd113,7'd14}:		p = 14'd1582;
            {7'd113,7'd15}:		p = 14'd1695;
            {7'd113,7'd16}:		p = 14'd1808;
            {7'd113,7'd17}:		p = 14'd1921;
            {7'd113,7'd18}:		p = 14'd2034;
            {7'd113,7'd19}:		p = 14'd2147;
            {7'd113,7'd20}:		p = 14'd2260;
            {7'd113,7'd21}:		p = 14'd2373;
            {7'd113,7'd22}:		p = 14'd2486;
            {7'd113,7'd23}:		p = 14'd2599;
            {7'd113,7'd24}:		p = 14'd2712;
            {7'd113,7'd25}:		p = 14'd2825;
            {7'd113,7'd26}:		p = 14'd2938;
            {7'd113,7'd27}:		p = 14'd3051;
            {7'd113,7'd28}:		p = 14'd3164;
            {7'd113,7'd29}:		p = 14'd3277;
            {7'd113,7'd30}:		p = 14'd3390;
            {7'd113,7'd31}:		p = 14'd3503;
            {7'd113,7'd32}:		p = 14'd3616;
            {7'd113,7'd33}:		p = 14'd3729;
            {7'd113,7'd34}:		p = 14'd3842;
            {7'd113,7'd35}:		p = 14'd3955;
            {7'd113,7'd36}:		p = 14'd4068;
            {7'd113,7'd37}:		p = 14'd4181;
            {7'd113,7'd38}:		p = 14'd4294;
            {7'd113,7'd39}:		p = 14'd4407;
            {7'd113,7'd40}:		p = 14'd4520;
            {7'd113,7'd41}:		p = 14'd4633;
            {7'd113,7'd42}:		p = 14'd4746;
            {7'd113,7'd43}:		p = 14'd4859;
            {7'd113,7'd44}:		p = 14'd4972;
            {7'd113,7'd45}:		p = 14'd5085;
            {7'd113,7'd46}:		p = 14'd5198;
            {7'd113,7'd47}:		p = 14'd5311;
            {7'd113,7'd48}:		p = 14'd5424;
            {7'd113,7'd49}:		p = 14'd5537;
            {7'd113,7'd50}:		p = 14'd5650;
            {7'd113,7'd51}:		p = 14'd5763;
            {7'd113,7'd52}:		p = 14'd5876;
            {7'd113,7'd53}:		p = 14'd5989;
            {7'd113,7'd54}:		p = 14'd6102;
            {7'd113,7'd55}:		p = 14'd6215;
            {7'd113,7'd56}:		p = 14'd6328;
            {7'd113,7'd57}:		p = 14'd6441;
            {7'd113,7'd58}:		p = 14'd6554;
            {7'd113,7'd59}:		p = 14'd6667;
            {7'd113,7'd60}:		p = 14'd6780;
            {7'd113,7'd61}:		p = 14'd6893;
            {7'd113,7'd62}:		p = 14'd7006;
            {7'd113,7'd63}:		p = 14'd7119;
            {7'd113,7'd64}:		p = 14'd7232;
            {7'd113,7'd65}:		p = 14'd7345;
            {7'd113,7'd66}:		p = 14'd7458;
            {7'd113,7'd67}:		p = 14'd7571;
            {7'd113,7'd68}:		p = 14'd7684;
            {7'd113,7'd69}:		p = 14'd7797;
            {7'd113,7'd70}:		p = 14'd7910;
            {7'd113,7'd71}:		p = 14'd8023;
            {7'd113,7'd72}:		p = 14'd8136;
            {7'd113,7'd73}:		p = 14'd8249;
            {7'd113,7'd74}:		p = 14'd8362;
            {7'd113,7'd75}:		p = 14'd8475;
            {7'd113,7'd76}:		p = 14'd8588;
            {7'd113,7'd77}:		p = 14'd8701;
            {7'd113,7'd78}:		p = 14'd8814;
            {7'd113,7'd79}:		p = 14'd8927;
            {7'd113,7'd80}:		p = 14'd9040;
            {7'd113,7'd81}:		p = 14'd9153;
            {7'd113,7'd82}:		p = 14'd9266;
            {7'd113,7'd83}:		p = 14'd9379;
            {7'd113,7'd84}:		p = 14'd9492;
            {7'd113,7'd85}:		p = 14'd9605;
            {7'd113,7'd86}:		p = 14'd9718;
            {7'd113,7'd87}:		p = 14'd9831;
            {7'd113,7'd88}:		p = 14'd9944;
            {7'd113,7'd89}:		p = 14'd10057;
            {7'd113,7'd90}:		p = 14'd10170;
            {7'd113,7'd91}:		p = 14'd10283;
            {7'd113,7'd92}:		p = 14'd10396;
            {7'd113,7'd93}:		p = 14'd10509;
            {7'd113,7'd94}:		p = 14'd10622;
            {7'd113,7'd95}:		p = 14'd10735;
            {7'd113,7'd96}:		p = 14'd10848;
            {7'd113,7'd97}:		p = 14'd10961;
            {7'd113,7'd98}:		p = 14'd11074;
            {7'd113,7'd99}:		p = 14'd11187;
            {7'd113,7'd100}:		p = 14'd11300;
            {7'd113,7'd101}:		p = 14'd11413;
            {7'd113,7'd102}:		p = 14'd11526;
            {7'd113,7'd103}:		p = 14'd11639;
            {7'd113,7'd104}:		p = 14'd11752;
            {7'd113,7'd105}:		p = 14'd11865;
            {7'd113,7'd106}:		p = 14'd11978;
            {7'd113,7'd107}:		p = 14'd12091;
            {7'd113,7'd108}:		p = 14'd12204;
            {7'd113,7'd109}:		p = 14'd12317;
            {7'd113,7'd110}:		p = 14'd12430;
            {7'd113,7'd111}:		p = 14'd12543;
            {7'd113,7'd112}:		p = 14'd12656;
            {7'd113,7'd113}:		p = 14'd12769;
            {7'd113,7'd114}:		p = 14'd12882;
            {7'd113,7'd115}:		p = 14'd12995;
            {7'd113,7'd116}:		p = 14'd13108;
            {7'd113,7'd117}:		p = 14'd13221;
            {7'd113,7'd118}:		p = 14'd13334;
            {7'd113,7'd119}:		p = 14'd13447;
            {7'd113,7'd120}:		p = 14'd13560;
            {7'd113,7'd121}:		p = 14'd13673;
            {7'd113,7'd122}:		p = 14'd13786;
            {7'd113,7'd123}:		p = 14'd13899;
            {7'd113,7'd124}:		p = 14'd14012;
            {7'd113,7'd125}:		p = 14'd14125;
            {7'd113,7'd126}:		p = 14'd14238;
            {7'd113,7'd127}:		p = 14'd14351;
            {7'd114,7'd0}:		p = 14'd0;
            {7'd114,7'd1}:		p = 14'd114;
            {7'd114,7'd2}:		p = 14'd228;
            {7'd114,7'd3}:		p = 14'd342;
            {7'd114,7'd4}:		p = 14'd456;
            {7'd114,7'd5}:		p = 14'd570;
            {7'd114,7'd6}:		p = 14'd684;
            {7'd114,7'd7}:		p = 14'd798;
            {7'd114,7'd8}:		p = 14'd912;
            {7'd114,7'd9}:		p = 14'd1026;
            {7'd114,7'd10}:		p = 14'd1140;
            {7'd114,7'd11}:		p = 14'd1254;
            {7'd114,7'd12}:		p = 14'd1368;
            {7'd114,7'd13}:		p = 14'd1482;
            {7'd114,7'd14}:		p = 14'd1596;
            {7'd114,7'd15}:		p = 14'd1710;
            {7'd114,7'd16}:		p = 14'd1824;
            {7'd114,7'd17}:		p = 14'd1938;
            {7'd114,7'd18}:		p = 14'd2052;
            {7'd114,7'd19}:		p = 14'd2166;
            {7'd114,7'd20}:		p = 14'd2280;
            {7'd114,7'd21}:		p = 14'd2394;
            {7'd114,7'd22}:		p = 14'd2508;
            {7'd114,7'd23}:		p = 14'd2622;
            {7'd114,7'd24}:		p = 14'd2736;
            {7'd114,7'd25}:		p = 14'd2850;
            {7'd114,7'd26}:		p = 14'd2964;
            {7'd114,7'd27}:		p = 14'd3078;
            {7'd114,7'd28}:		p = 14'd3192;
            {7'd114,7'd29}:		p = 14'd3306;
            {7'd114,7'd30}:		p = 14'd3420;
            {7'd114,7'd31}:		p = 14'd3534;
            {7'd114,7'd32}:		p = 14'd3648;
            {7'd114,7'd33}:		p = 14'd3762;
            {7'd114,7'd34}:		p = 14'd3876;
            {7'd114,7'd35}:		p = 14'd3990;
            {7'd114,7'd36}:		p = 14'd4104;
            {7'd114,7'd37}:		p = 14'd4218;
            {7'd114,7'd38}:		p = 14'd4332;
            {7'd114,7'd39}:		p = 14'd4446;
            {7'd114,7'd40}:		p = 14'd4560;
            {7'd114,7'd41}:		p = 14'd4674;
            {7'd114,7'd42}:		p = 14'd4788;
            {7'd114,7'd43}:		p = 14'd4902;
            {7'd114,7'd44}:		p = 14'd5016;
            {7'd114,7'd45}:		p = 14'd5130;
            {7'd114,7'd46}:		p = 14'd5244;
            {7'd114,7'd47}:		p = 14'd5358;
            {7'd114,7'd48}:		p = 14'd5472;
            {7'd114,7'd49}:		p = 14'd5586;
            {7'd114,7'd50}:		p = 14'd5700;
            {7'd114,7'd51}:		p = 14'd5814;
            {7'd114,7'd52}:		p = 14'd5928;
            {7'd114,7'd53}:		p = 14'd6042;
            {7'd114,7'd54}:		p = 14'd6156;
            {7'd114,7'd55}:		p = 14'd6270;
            {7'd114,7'd56}:		p = 14'd6384;
            {7'd114,7'd57}:		p = 14'd6498;
            {7'd114,7'd58}:		p = 14'd6612;
            {7'd114,7'd59}:		p = 14'd6726;
            {7'd114,7'd60}:		p = 14'd6840;
            {7'd114,7'd61}:		p = 14'd6954;
            {7'd114,7'd62}:		p = 14'd7068;
            {7'd114,7'd63}:		p = 14'd7182;
            {7'd114,7'd64}:		p = 14'd7296;
            {7'd114,7'd65}:		p = 14'd7410;
            {7'd114,7'd66}:		p = 14'd7524;
            {7'd114,7'd67}:		p = 14'd7638;
            {7'd114,7'd68}:		p = 14'd7752;
            {7'd114,7'd69}:		p = 14'd7866;
            {7'd114,7'd70}:		p = 14'd7980;
            {7'd114,7'd71}:		p = 14'd8094;
            {7'd114,7'd72}:		p = 14'd8208;
            {7'd114,7'd73}:		p = 14'd8322;
            {7'd114,7'd74}:		p = 14'd8436;
            {7'd114,7'd75}:		p = 14'd8550;
            {7'd114,7'd76}:		p = 14'd8664;
            {7'd114,7'd77}:		p = 14'd8778;
            {7'd114,7'd78}:		p = 14'd8892;
            {7'd114,7'd79}:		p = 14'd9006;
            {7'd114,7'd80}:		p = 14'd9120;
            {7'd114,7'd81}:		p = 14'd9234;
            {7'd114,7'd82}:		p = 14'd9348;
            {7'd114,7'd83}:		p = 14'd9462;
            {7'd114,7'd84}:		p = 14'd9576;
            {7'd114,7'd85}:		p = 14'd9690;
            {7'd114,7'd86}:		p = 14'd9804;
            {7'd114,7'd87}:		p = 14'd9918;
            {7'd114,7'd88}:		p = 14'd10032;
            {7'd114,7'd89}:		p = 14'd10146;
            {7'd114,7'd90}:		p = 14'd10260;
            {7'd114,7'd91}:		p = 14'd10374;
            {7'd114,7'd92}:		p = 14'd10488;
            {7'd114,7'd93}:		p = 14'd10602;
            {7'd114,7'd94}:		p = 14'd10716;
            {7'd114,7'd95}:		p = 14'd10830;
            {7'd114,7'd96}:		p = 14'd10944;
            {7'd114,7'd97}:		p = 14'd11058;
            {7'd114,7'd98}:		p = 14'd11172;
            {7'd114,7'd99}:		p = 14'd11286;
            {7'd114,7'd100}:		p = 14'd11400;
            {7'd114,7'd101}:		p = 14'd11514;
            {7'd114,7'd102}:		p = 14'd11628;
            {7'd114,7'd103}:		p = 14'd11742;
            {7'd114,7'd104}:		p = 14'd11856;
            {7'd114,7'd105}:		p = 14'd11970;
            {7'd114,7'd106}:		p = 14'd12084;
            {7'd114,7'd107}:		p = 14'd12198;
            {7'd114,7'd108}:		p = 14'd12312;
            {7'd114,7'd109}:		p = 14'd12426;
            {7'd114,7'd110}:		p = 14'd12540;
            {7'd114,7'd111}:		p = 14'd12654;
            {7'd114,7'd112}:		p = 14'd12768;
            {7'd114,7'd113}:		p = 14'd12882;
            {7'd114,7'd114}:		p = 14'd12996;
            {7'd114,7'd115}:		p = 14'd13110;
            {7'd114,7'd116}:		p = 14'd13224;
            {7'd114,7'd117}:		p = 14'd13338;
            {7'd114,7'd118}:		p = 14'd13452;
            {7'd114,7'd119}:		p = 14'd13566;
            {7'd114,7'd120}:		p = 14'd13680;
            {7'd114,7'd121}:		p = 14'd13794;
            {7'd114,7'd122}:		p = 14'd13908;
            {7'd114,7'd123}:		p = 14'd14022;
            {7'd114,7'd124}:		p = 14'd14136;
            {7'd114,7'd125}:		p = 14'd14250;
            {7'd114,7'd126}:		p = 14'd14364;
            {7'd114,7'd127}:		p = 14'd14478;
            {7'd115,7'd0}:		p = 14'd0;
            {7'd115,7'd1}:		p = 14'd115;
            {7'd115,7'd2}:		p = 14'd230;
            {7'd115,7'd3}:		p = 14'd345;
            {7'd115,7'd4}:		p = 14'd460;
            {7'd115,7'd5}:		p = 14'd575;
            {7'd115,7'd6}:		p = 14'd690;
            {7'd115,7'd7}:		p = 14'd805;
            {7'd115,7'd8}:		p = 14'd920;
            {7'd115,7'd9}:		p = 14'd1035;
            {7'd115,7'd10}:		p = 14'd1150;
            {7'd115,7'd11}:		p = 14'd1265;
            {7'd115,7'd12}:		p = 14'd1380;
            {7'd115,7'd13}:		p = 14'd1495;
            {7'd115,7'd14}:		p = 14'd1610;
            {7'd115,7'd15}:		p = 14'd1725;
            {7'd115,7'd16}:		p = 14'd1840;
            {7'd115,7'd17}:		p = 14'd1955;
            {7'd115,7'd18}:		p = 14'd2070;
            {7'd115,7'd19}:		p = 14'd2185;
            {7'd115,7'd20}:		p = 14'd2300;
            {7'd115,7'd21}:		p = 14'd2415;
            {7'd115,7'd22}:		p = 14'd2530;
            {7'd115,7'd23}:		p = 14'd2645;
            {7'd115,7'd24}:		p = 14'd2760;
            {7'd115,7'd25}:		p = 14'd2875;
            {7'd115,7'd26}:		p = 14'd2990;
            {7'd115,7'd27}:		p = 14'd3105;
            {7'd115,7'd28}:		p = 14'd3220;
            {7'd115,7'd29}:		p = 14'd3335;
            {7'd115,7'd30}:		p = 14'd3450;
            {7'd115,7'd31}:		p = 14'd3565;
            {7'd115,7'd32}:		p = 14'd3680;
            {7'd115,7'd33}:		p = 14'd3795;
            {7'd115,7'd34}:		p = 14'd3910;
            {7'd115,7'd35}:		p = 14'd4025;
            {7'd115,7'd36}:		p = 14'd4140;
            {7'd115,7'd37}:		p = 14'd4255;
            {7'd115,7'd38}:		p = 14'd4370;
            {7'd115,7'd39}:		p = 14'd4485;
            {7'd115,7'd40}:		p = 14'd4600;
            {7'd115,7'd41}:		p = 14'd4715;
            {7'd115,7'd42}:		p = 14'd4830;
            {7'd115,7'd43}:		p = 14'd4945;
            {7'd115,7'd44}:		p = 14'd5060;
            {7'd115,7'd45}:		p = 14'd5175;
            {7'd115,7'd46}:		p = 14'd5290;
            {7'd115,7'd47}:		p = 14'd5405;
            {7'd115,7'd48}:		p = 14'd5520;
            {7'd115,7'd49}:		p = 14'd5635;
            {7'd115,7'd50}:		p = 14'd5750;
            {7'd115,7'd51}:		p = 14'd5865;
            {7'd115,7'd52}:		p = 14'd5980;
            {7'd115,7'd53}:		p = 14'd6095;
            {7'd115,7'd54}:		p = 14'd6210;
            {7'd115,7'd55}:		p = 14'd6325;
            {7'd115,7'd56}:		p = 14'd6440;
            {7'd115,7'd57}:		p = 14'd6555;
            {7'd115,7'd58}:		p = 14'd6670;
            {7'd115,7'd59}:		p = 14'd6785;
            {7'd115,7'd60}:		p = 14'd6900;
            {7'd115,7'd61}:		p = 14'd7015;
            {7'd115,7'd62}:		p = 14'd7130;
            {7'd115,7'd63}:		p = 14'd7245;
            {7'd115,7'd64}:		p = 14'd7360;
            {7'd115,7'd65}:		p = 14'd7475;
            {7'd115,7'd66}:		p = 14'd7590;
            {7'd115,7'd67}:		p = 14'd7705;
            {7'd115,7'd68}:		p = 14'd7820;
            {7'd115,7'd69}:		p = 14'd7935;
            {7'd115,7'd70}:		p = 14'd8050;
            {7'd115,7'd71}:		p = 14'd8165;
            {7'd115,7'd72}:		p = 14'd8280;
            {7'd115,7'd73}:		p = 14'd8395;
            {7'd115,7'd74}:		p = 14'd8510;
            {7'd115,7'd75}:		p = 14'd8625;
            {7'd115,7'd76}:		p = 14'd8740;
            {7'd115,7'd77}:		p = 14'd8855;
            {7'd115,7'd78}:		p = 14'd8970;
            {7'd115,7'd79}:		p = 14'd9085;
            {7'd115,7'd80}:		p = 14'd9200;
            {7'd115,7'd81}:		p = 14'd9315;
            {7'd115,7'd82}:		p = 14'd9430;
            {7'd115,7'd83}:		p = 14'd9545;
            {7'd115,7'd84}:		p = 14'd9660;
            {7'd115,7'd85}:		p = 14'd9775;
            {7'd115,7'd86}:		p = 14'd9890;
            {7'd115,7'd87}:		p = 14'd10005;
            {7'd115,7'd88}:		p = 14'd10120;
            {7'd115,7'd89}:		p = 14'd10235;
            {7'd115,7'd90}:		p = 14'd10350;
            {7'd115,7'd91}:		p = 14'd10465;
            {7'd115,7'd92}:		p = 14'd10580;
            {7'd115,7'd93}:		p = 14'd10695;
            {7'd115,7'd94}:		p = 14'd10810;
            {7'd115,7'd95}:		p = 14'd10925;
            {7'd115,7'd96}:		p = 14'd11040;
            {7'd115,7'd97}:		p = 14'd11155;
            {7'd115,7'd98}:		p = 14'd11270;
            {7'd115,7'd99}:		p = 14'd11385;
            {7'd115,7'd100}:		p = 14'd11500;
            {7'd115,7'd101}:		p = 14'd11615;
            {7'd115,7'd102}:		p = 14'd11730;
            {7'd115,7'd103}:		p = 14'd11845;
            {7'd115,7'd104}:		p = 14'd11960;
            {7'd115,7'd105}:		p = 14'd12075;
            {7'd115,7'd106}:		p = 14'd12190;
            {7'd115,7'd107}:		p = 14'd12305;
            {7'd115,7'd108}:		p = 14'd12420;
            {7'd115,7'd109}:		p = 14'd12535;
            {7'd115,7'd110}:		p = 14'd12650;
            {7'd115,7'd111}:		p = 14'd12765;
            {7'd115,7'd112}:		p = 14'd12880;
            {7'd115,7'd113}:		p = 14'd12995;
            {7'd115,7'd114}:		p = 14'd13110;
            {7'd115,7'd115}:		p = 14'd13225;
            {7'd115,7'd116}:		p = 14'd13340;
            {7'd115,7'd117}:		p = 14'd13455;
            {7'd115,7'd118}:		p = 14'd13570;
            {7'd115,7'd119}:		p = 14'd13685;
            {7'd115,7'd120}:		p = 14'd13800;
            {7'd115,7'd121}:		p = 14'd13915;
            {7'd115,7'd122}:		p = 14'd14030;
            {7'd115,7'd123}:		p = 14'd14145;
            {7'd115,7'd124}:		p = 14'd14260;
            {7'd115,7'd125}:		p = 14'd14375;
            {7'd115,7'd126}:		p = 14'd14490;
            {7'd115,7'd127}:		p = 14'd14605;
            {7'd116,7'd0}:		p = 14'd0;
            {7'd116,7'd1}:		p = 14'd116;
            {7'd116,7'd2}:		p = 14'd232;
            {7'd116,7'd3}:		p = 14'd348;
            {7'd116,7'd4}:		p = 14'd464;
            {7'd116,7'd5}:		p = 14'd580;
            {7'd116,7'd6}:		p = 14'd696;
            {7'd116,7'd7}:		p = 14'd812;
            {7'd116,7'd8}:		p = 14'd928;
            {7'd116,7'd9}:		p = 14'd1044;
            {7'd116,7'd10}:		p = 14'd1160;
            {7'd116,7'd11}:		p = 14'd1276;
            {7'd116,7'd12}:		p = 14'd1392;
            {7'd116,7'd13}:		p = 14'd1508;
            {7'd116,7'd14}:		p = 14'd1624;
            {7'd116,7'd15}:		p = 14'd1740;
            {7'd116,7'd16}:		p = 14'd1856;
            {7'd116,7'd17}:		p = 14'd1972;
            {7'd116,7'd18}:		p = 14'd2088;
            {7'd116,7'd19}:		p = 14'd2204;
            {7'd116,7'd20}:		p = 14'd2320;
            {7'd116,7'd21}:		p = 14'd2436;
            {7'd116,7'd22}:		p = 14'd2552;
            {7'd116,7'd23}:		p = 14'd2668;
            {7'd116,7'd24}:		p = 14'd2784;
            {7'd116,7'd25}:		p = 14'd2900;
            {7'd116,7'd26}:		p = 14'd3016;
            {7'd116,7'd27}:		p = 14'd3132;
            {7'd116,7'd28}:		p = 14'd3248;
            {7'd116,7'd29}:		p = 14'd3364;
            {7'd116,7'd30}:		p = 14'd3480;
            {7'd116,7'd31}:		p = 14'd3596;
            {7'd116,7'd32}:		p = 14'd3712;
            {7'd116,7'd33}:		p = 14'd3828;
            {7'd116,7'd34}:		p = 14'd3944;
            {7'd116,7'd35}:		p = 14'd4060;
            {7'd116,7'd36}:		p = 14'd4176;
            {7'd116,7'd37}:		p = 14'd4292;
            {7'd116,7'd38}:		p = 14'd4408;
            {7'd116,7'd39}:		p = 14'd4524;
            {7'd116,7'd40}:		p = 14'd4640;
            {7'd116,7'd41}:		p = 14'd4756;
            {7'd116,7'd42}:		p = 14'd4872;
            {7'd116,7'd43}:		p = 14'd4988;
            {7'd116,7'd44}:		p = 14'd5104;
            {7'd116,7'd45}:		p = 14'd5220;
            {7'd116,7'd46}:		p = 14'd5336;
            {7'd116,7'd47}:		p = 14'd5452;
            {7'd116,7'd48}:		p = 14'd5568;
            {7'd116,7'd49}:		p = 14'd5684;
            {7'd116,7'd50}:		p = 14'd5800;
            {7'd116,7'd51}:		p = 14'd5916;
            {7'd116,7'd52}:		p = 14'd6032;
            {7'd116,7'd53}:		p = 14'd6148;
            {7'd116,7'd54}:		p = 14'd6264;
            {7'd116,7'd55}:		p = 14'd6380;
            {7'd116,7'd56}:		p = 14'd6496;
            {7'd116,7'd57}:		p = 14'd6612;
            {7'd116,7'd58}:		p = 14'd6728;
            {7'd116,7'd59}:		p = 14'd6844;
            {7'd116,7'd60}:		p = 14'd6960;
            {7'd116,7'd61}:		p = 14'd7076;
            {7'd116,7'd62}:		p = 14'd7192;
            {7'd116,7'd63}:		p = 14'd7308;
            {7'd116,7'd64}:		p = 14'd7424;
            {7'd116,7'd65}:		p = 14'd7540;
            {7'd116,7'd66}:		p = 14'd7656;
            {7'd116,7'd67}:		p = 14'd7772;
            {7'd116,7'd68}:		p = 14'd7888;
            {7'd116,7'd69}:		p = 14'd8004;
            {7'd116,7'd70}:		p = 14'd8120;
            {7'd116,7'd71}:		p = 14'd8236;
            {7'd116,7'd72}:		p = 14'd8352;
            {7'd116,7'd73}:		p = 14'd8468;
            {7'd116,7'd74}:		p = 14'd8584;
            {7'd116,7'd75}:		p = 14'd8700;
            {7'd116,7'd76}:		p = 14'd8816;
            {7'd116,7'd77}:		p = 14'd8932;
            {7'd116,7'd78}:		p = 14'd9048;
            {7'd116,7'd79}:		p = 14'd9164;
            {7'd116,7'd80}:		p = 14'd9280;
            {7'd116,7'd81}:		p = 14'd9396;
            {7'd116,7'd82}:		p = 14'd9512;
            {7'd116,7'd83}:		p = 14'd9628;
            {7'd116,7'd84}:		p = 14'd9744;
            {7'd116,7'd85}:		p = 14'd9860;
            {7'd116,7'd86}:		p = 14'd9976;
            {7'd116,7'd87}:		p = 14'd10092;
            {7'd116,7'd88}:		p = 14'd10208;
            {7'd116,7'd89}:		p = 14'd10324;
            {7'd116,7'd90}:		p = 14'd10440;
            {7'd116,7'd91}:		p = 14'd10556;
            {7'd116,7'd92}:		p = 14'd10672;
            {7'd116,7'd93}:		p = 14'd10788;
            {7'd116,7'd94}:		p = 14'd10904;
            {7'd116,7'd95}:		p = 14'd11020;
            {7'd116,7'd96}:		p = 14'd11136;
            {7'd116,7'd97}:		p = 14'd11252;
            {7'd116,7'd98}:		p = 14'd11368;
            {7'd116,7'd99}:		p = 14'd11484;
            {7'd116,7'd100}:		p = 14'd11600;
            {7'd116,7'd101}:		p = 14'd11716;
            {7'd116,7'd102}:		p = 14'd11832;
            {7'd116,7'd103}:		p = 14'd11948;
            {7'd116,7'd104}:		p = 14'd12064;
            {7'd116,7'd105}:		p = 14'd12180;
            {7'd116,7'd106}:		p = 14'd12296;
            {7'd116,7'd107}:		p = 14'd12412;
            {7'd116,7'd108}:		p = 14'd12528;
            {7'd116,7'd109}:		p = 14'd12644;
            {7'd116,7'd110}:		p = 14'd12760;
            {7'd116,7'd111}:		p = 14'd12876;
            {7'd116,7'd112}:		p = 14'd12992;
            {7'd116,7'd113}:		p = 14'd13108;
            {7'd116,7'd114}:		p = 14'd13224;
            {7'd116,7'd115}:		p = 14'd13340;
            {7'd116,7'd116}:		p = 14'd13456;
            {7'd116,7'd117}:		p = 14'd13572;
            {7'd116,7'd118}:		p = 14'd13688;
            {7'd116,7'd119}:		p = 14'd13804;
            {7'd116,7'd120}:		p = 14'd13920;
            {7'd116,7'd121}:		p = 14'd14036;
            {7'd116,7'd122}:		p = 14'd14152;
            {7'd116,7'd123}:		p = 14'd14268;
            {7'd116,7'd124}:		p = 14'd14384;
            {7'd116,7'd125}:		p = 14'd14500;
            {7'd116,7'd126}:		p = 14'd14616;
            {7'd116,7'd127}:		p = 14'd14732;
            {7'd117,7'd0}:		p = 14'd0;
            {7'd117,7'd1}:		p = 14'd117;
            {7'd117,7'd2}:		p = 14'd234;
            {7'd117,7'd3}:		p = 14'd351;
            {7'd117,7'd4}:		p = 14'd468;
            {7'd117,7'd5}:		p = 14'd585;
            {7'd117,7'd6}:		p = 14'd702;
            {7'd117,7'd7}:		p = 14'd819;
            {7'd117,7'd8}:		p = 14'd936;
            {7'd117,7'd9}:		p = 14'd1053;
            {7'd117,7'd10}:		p = 14'd1170;
            {7'd117,7'd11}:		p = 14'd1287;
            {7'd117,7'd12}:		p = 14'd1404;
            {7'd117,7'd13}:		p = 14'd1521;
            {7'd117,7'd14}:		p = 14'd1638;
            {7'd117,7'd15}:		p = 14'd1755;
            {7'd117,7'd16}:		p = 14'd1872;
            {7'd117,7'd17}:		p = 14'd1989;
            {7'd117,7'd18}:		p = 14'd2106;
            {7'd117,7'd19}:		p = 14'd2223;
            {7'd117,7'd20}:		p = 14'd2340;
            {7'd117,7'd21}:		p = 14'd2457;
            {7'd117,7'd22}:		p = 14'd2574;
            {7'd117,7'd23}:		p = 14'd2691;
            {7'd117,7'd24}:		p = 14'd2808;
            {7'd117,7'd25}:		p = 14'd2925;
            {7'd117,7'd26}:		p = 14'd3042;
            {7'd117,7'd27}:		p = 14'd3159;
            {7'd117,7'd28}:		p = 14'd3276;
            {7'd117,7'd29}:		p = 14'd3393;
            {7'd117,7'd30}:		p = 14'd3510;
            {7'd117,7'd31}:		p = 14'd3627;
            {7'd117,7'd32}:		p = 14'd3744;
            {7'd117,7'd33}:		p = 14'd3861;
            {7'd117,7'd34}:		p = 14'd3978;
            {7'd117,7'd35}:		p = 14'd4095;
            {7'd117,7'd36}:		p = 14'd4212;
            {7'd117,7'd37}:		p = 14'd4329;
            {7'd117,7'd38}:		p = 14'd4446;
            {7'd117,7'd39}:		p = 14'd4563;
            {7'd117,7'd40}:		p = 14'd4680;
            {7'd117,7'd41}:		p = 14'd4797;
            {7'd117,7'd42}:		p = 14'd4914;
            {7'd117,7'd43}:		p = 14'd5031;
            {7'd117,7'd44}:		p = 14'd5148;
            {7'd117,7'd45}:		p = 14'd5265;
            {7'd117,7'd46}:		p = 14'd5382;
            {7'd117,7'd47}:		p = 14'd5499;
            {7'd117,7'd48}:		p = 14'd5616;
            {7'd117,7'd49}:		p = 14'd5733;
            {7'd117,7'd50}:		p = 14'd5850;
            {7'd117,7'd51}:		p = 14'd5967;
            {7'd117,7'd52}:		p = 14'd6084;
            {7'd117,7'd53}:		p = 14'd6201;
            {7'd117,7'd54}:		p = 14'd6318;
            {7'd117,7'd55}:		p = 14'd6435;
            {7'd117,7'd56}:		p = 14'd6552;
            {7'd117,7'd57}:		p = 14'd6669;
            {7'd117,7'd58}:		p = 14'd6786;
            {7'd117,7'd59}:		p = 14'd6903;
            {7'd117,7'd60}:		p = 14'd7020;
            {7'd117,7'd61}:		p = 14'd7137;
            {7'd117,7'd62}:		p = 14'd7254;
            {7'd117,7'd63}:		p = 14'd7371;
            {7'd117,7'd64}:		p = 14'd7488;
            {7'd117,7'd65}:		p = 14'd7605;
            {7'd117,7'd66}:		p = 14'd7722;
            {7'd117,7'd67}:		p = 14'd7839;
            {7'd117,7'd68}:		p = 14'd7956;
            {7'd117,7'd69}:		p = 14'd8073;
            {7'd117,7'd70}:		p = 14'd8190;
            {7'd117,7'd71}:		p = 14'd8307;
            {7'd117,7'd72}:		p = 14'd8424;
            {7'd117,7'd73}:		p = 14'd8541;
            {7'd117,7'd74}:		p = 14'd8658;
            {7'd117,7'd75}:		p = 14'd8775;
            {7'd117,7'd76}:		p = 14'd8892;
            {7'd117,7'd77}:		p = 14'd9009;
            {7'd117,7'd78}:		p = 14'd9126;
            {7'd117,7'd79}:		p = 14'd9243;
            {7'd117,7'd80}:		p = 14'd9360;
            {7'd117,7'd81}:		p = 14'd9477;
            {7'd117,7'd82}:		p = 14'd9594;
            {7'd117,7'd83}:		p = 14'd9711;
            {7'd117,7'd84}:		p = 14'd9828;
            {7'd117,7'd85}:		p = 14'd9945;
            {7'd117,7'd86}:		p = 14'd10062;
            {7'd117,7'd87}:		p = 14'd10179;
            {7'd117,7'd88}:		p = 14'd10296;
            {7'd117,7'd89}:		p = 14'd10413;
            {7'd117,7'd90}:		p = 14'd10530;
            {7'd117,7'd91}:		p = 14'd10647;
            {7'd117,7'd92}:		p = 14'd10764;
            {7'd117,7'd93}:		p = 14'd10881;
            {7'd117,7'd94}:		p = 14'd10998;
            {7'd117,7'd95}:		p = 14'd11115;
            {7'd117,7'd96}:		p = 14'd11232;
            {7'd117,7'd97}:		p = 14'd11349;
            {7'd117,7'd98}:		p = 14'd11466;
            {7'd117,7'd99}:		p = 14'd11583;
            {7'd117,7'd100}:		p = 14'd11700;
            {7'd117,7'd101}:		p = 14'd11817;
            {7'd117,7'd102}:		p = 14'd11934;
            {7'd117,7'd103}:		p = 14'd12051;
            {7'd117,7'd104}:		p = 14'd12168;
            {7'd117,7'd105}:		p = 14'd12285;
            {7'd117,7'd106}:		p = 14'd12402;
            {7'd117,7'd107}:		p = 14'd12519;
            {7'd117,7'd108}:		p = 14'd12636;
            {7'd117,7'd109}:		p = 14'd12753;
            {7'd117,7'd110}:		p = 14'd12870;
            {7'd117,7'd111}:		p = 14'd12987;
            {7'd117,7'd112}:		p = 14'd13104;
            {7'd117,7'd113}:		p = 14'd13221;
            {7'd117,7'd114}:		p = 14'd13338;
            {7'd117,7'd115}:		p = 14'd13455;
            {7'd117,7'd116}:		p = 14'd13572;
            {7'd117,7'd117}:		p = 14'd13689;
            {7'd117,7'd118}:		p = 14'd13806;
            {7'd117,7'd119}:		p = 14'd13923;
            {7'd117,7'd120}:		p = 14'd14040;
            {7'd117,7'd121}:		p = 14'd14157;
            {7'd117,7'd122}:		p = 14'd14274;
            {7'd117,7'd123}:		p = 14'd14391;
            {7'd117,7'd124}:		p = 14'd14508;
            {7'd117,7'd125}:		p = 14'd14625;
            {7'd117,7'd126}:		p = 14'd14742;
            {7'd117,7'd127}:		p = 14'd14859;
            {7'd118,7'd0}:		p = 14'd0;
            {7'd118,7'd1}:		p = 14'd118;
            {7'd118,7'd2}:		p = 14'd236;
            {7'd118,7'd3}:		p = 14'd354;
            {7'd118,7'd4}:		p = 14'd472;
            {7'd118,7'd5}:		p = 14'd590;
            {7'd118,7'd6}:		p = 14'd708;
            {7'd118,7'd7}:		p = 14'd826;
            {7'd118,7'd8}:		p = 14'd944;
            {7'd118,7'd9}:		p = 14'd1062;
            {7'd118,7'd10}:		p = 14'd1180;
            {7'd118,7'd11}:		p = 14'd1298;
            {7'd118,7'd12}:		p = 14'd1416;
            {7'd118,7'd13}:		p = 14'd1534;
            {7'd118,7'd14}:		p = 14'd1652;
            {7'd118,7'd15}:		p = 14'd1770;
            {7'd118,7'd16}:		p = 14'd1888;
            {7'd118,7'd17}:		p = 14'd2006;
            {7'd118,7'd18}:		p = 14'd2124;
            {7'd118,7'd19}:		p = 14'd2242;
            {7'd118,7'd20}:		p = 14'd2360;
            {7'd118,7'd21}:		p = 14'd2478;
            {7'd118,7'd22}:		p = 14'd2596;
            {7'd118,7'd23}:		p = 14'd2714;
            {7'd118,7'd24}:		p = 14'd2832;
            {7'd118,7'd25}:		p = 14'd2950;
            {7'd118,7'd26}:		p = 14'd3068;
            {7'd118,7'd27}:		p = 14'd3186;
            {7'd118,7'd28}:		p = 14'd3304;
            {7'd118,7'd29}:		p = 14'd3422;
            {7'd118,7'd30}:		p = 14'd3540;
            {7'd118,7'd31}:		p = 14'd3658;
            {7'd118,7'd32}:		p = 14'd3776;
            {7'd118,7'd33}:		p = 14'd3894;
            {7'd118,7'd34}:		p = 14'd4012;
            {7'd118,7'd35}:		p = 14'd4130;
            {7'd118,7'd36}:		p = 14'd4248;
            {7'd118,7'd37}:		p = 14'd4366;
            {7'd118,7'd38}:		p = 14'd4484;
            {7'd118,7'd39}:		p = 14'd4602;
            {7'd118,7'd40}:		p = 14'd4720;
            {7'd118,7'd41}:		p = 14'd4838;
            {7'd118,7'd42}:		p = 14'd4956;
            {7'd118,7'd43}:		p = 14'd5074;
            {7'd118,7'd44}:		p = 14'd5192;
            {7'd118,7'd45}:		p = 14'd5310;
            {7'd118,7'd46}:		p = 14'd5428;
            {7'd118,7'd47}:		p = 14'd5546;
            {7'd118,7'd48}:		p = 14'd5664;
            {7'd118,7'd49}:		p = 14'd5782;
            {7'd118,7'd50}:		p = 14'd5900;
            {7'd118,7'd51}:		p = 14'd6018;
            {7'd118,7'd52}:		p = 14'd6136;
            {7'd118,7'd53}:		p = 14'd6254;
            {7'd118,7'd54}:		p = 14'd6372;
            {7'd118,7'd55}:		p = 14'd6490;
            {7'd118,7'd56}:		p = 14'd6608;
            {7'd118,7'd57}:		p = 14'd6726;
            {7'd118,7'd58}:		p = 14'd6844;
            {7'd118,7'd59}:		p = 14'd6962;
            {7'd118,7'd60}:		p = 14'd7080;
            {7'd118,7'd61}:		p = 14'd7198;
            {7'd118,7'd62}:		p = 14'd7316;
            {7'd118,7'd63}:		p = 14'd7434;
            {7'd118,7'd64}:		p = 14'd7552;
            {7'd118,7'd65}:		p = 14'd7670;
            {7'd118,7'd66}:		p = 14'd7788;
            {7'd118,7'd67}:		p = 14'd7906;
            {7'd118,7'd68}:		p = 14'd8024;
            {7'd118,7'd69}:		p = 14'd8142;
            {7'd118,7'd70}:		p = 14'd8260;
            {7'd118,7'd71}:		p = 14'd8378;
            {7'd118,7'd72}:		p = 14'd8496;
            {7'd118,7'd73}:		p = 14'd8614;
            {7'd118,7'd74}:		p = 14'd8732;
            {7'd118,7'd75}:		p = 14'd8850;
            {7'd118,7'd76}:		p = 14'd8968;
            {7'd118,7'd77}:		p = 14'd9086;
            {7'd118,7'd78}:		p = 14'd9204;
            {7'd118,7'd79}:		p = 14'd9322;
            {7'd118,7'd80}:		p = 14'd9440;
            {7'd118,7'd81}:		p = 14'd9558;
            {7'd118,7'd82}:		p = 14'd9676;
            {7'd118,7'd83}:		p = 14'd9794;
            {7'd118,7'd84}:		p = 14'd9912;
            {7'd118,7'd85}:		p = 14'd10030;
            {7'd118,7'd86}:		p = 14'd10148;
            {7'd118,7'd87}:		p = 14'd10266;
            {7'd118,7'd88}:		p = 14'd10384;
            {7'd118,7'd89}:		p = 14'd10502;
            {7'd118,7'd90}:		p = 14'd10620;
            {7'd118,7'd91}:		p = 14'd10738;
            {7'd118,7'd92}:		p = 14'd10856;
            {7'd118,7'd93}:		p = 14'd10974;
            {7'd118,7'd94}:		p = 14'd11092;
            {7'd118,7'd95}:		p = 14'd11210;
            {7'd118,7'd96}:		p = 14'd11328;
            {7'd118,7'd97}:		p = 14'd11446;
            {7'd118,7'd98}:		p = 14'd11564;
            {7'd118,7'd99}:		p = 14'd11682;
            {7'd118,7'd100}:		p = 14'd11800;
            {7'd118,7'd101}:		p = 14'd11918;
            {7'd118,7'd102}:		p = 14'd12036;
            {7'd118,7'd103}:		p = 14'd12154;
            {7'd118,7'd104}:		p = 14'd12272;
            {7'd118,7'd105}:		p = 14'd12390;
            {7'd118,7'd106}:		p = 14'd12508;
            {7'd118,7'd107}:		p = 14'd12626;
            {7'd118,7'd108}:		p = 14'd12744;
            {7'd118,7'd109}:		p = 14'd12862;
            {7'd118,7'd110}:		p = 14'd12980;
            {7'd118,7'd111}:		p = 14'd13098;
            {7'd118,7'd112}:		p = 14'd13216;
            {7'd118,7'd113}:		p = 14'd13334;
            {7'd118,7'd114}:		p = 14'd13452;
            {7'd118,7'd115}:		p = 14'd13570;
            {7'd118,7'd116}:		p = 14'd13688;
            {7'd118,7'd117}:		p = 14'd13806;
            {7'd118,7'd118}:		p = 14'd13924;
            {7'd118,7'd119}:		p = 14'd14042;
            {7'd118,7'd120}:		p = 14'd14160;
            {7'd118,7'd121}:		p = 14'd14278;
            {7'd118,7'd122}:		p = 14'd14396;
            {7'd118,7'd123}:		p = 14'd14514;
            {7'd118,7'd124}:		p = 14'd14632;
            {7'd118,7'd125}:		p = 14'd14750;
            {7'd118,7'd126}:		p = 14'd14868;
            {7'd118,7'd127}:		p = 14'd14986;
            {7'd119,7'd0}:		p = 14'd0;
            {7'd119,7'd1}:		p = 14'd119;
            {7'd119,7'd2}:		p = 14'd238;
            {7'd119,7'd3}:		p = 14'd357;
            {7'd119,7'd4}:		p = 14'd476;
            {7'd119,7'd5}:		p = 14'd595;
            {7'd119,7'd6}:		p = 14'd714;
            {7'd119,7'd7}:		p = 14'd833;
            {7'd119,7'd8}:		p = 14'd952;
            {7'd119,7'd9}:		p = 14'd1071;
            {7'd119,7'd10}:		p = 14'd1190;
            {7'd119,7'd11}:		p = 14'd1309;
            {7'd119,7'd12}:		p = 14'd1428;
            {7'd119,7'd13}:		p = 14'd1547;
            {7'd119,7'd14}:		p = 14'd1666;
            {7'd119,7'd15}:		p = 14'd1785;
            {7'd119,7'd16}:		p = 14'd1904;
            {7'd119,7'd17}:		p = 14'd2023;
            {7'd119,7'd18}:		p = 14'd2142;
            {7'd119,7'd19}:		p = 14'd2261;
            {7'd119,7'd20}:		p = 14'd2380;
            {7'd119,7'd21}:		p = 14'd2499;
            {7'd119,7'd22}:		p = 14'd2618;
            {7'd119,7'd23}:		p = 14'd2737;
            {7'd119,7'd24}:		p = 14'd2856;
            {7'd119,7'd25}:		p = 14'd2975;
            {7'd119,7'd26}:		p = 14'd3094;
            {7'd119,7'd27}:		p = 14'd3213;
            {7'd119,7'd28}:		p = 14'd3332;
            {7'd119,7'd29}:		p = 14'd3451;
            {7'd119,7'd30}:		p = 14'd3570;
            {7'd119,7'd31}:		p = 14'd3689;
            {7'd119,7'd32}:		p = 14'd3808;
            {7'd119,7'd33}:		p = 14'd3927;
            {7'd119,7'd34}:		p = 14'd4046;
            {7'd119,7'd35}:		p = 14'd4165;
            {7'd119,7'd36}:		p = 14'd4284;
            {7'd119,7'd37}:		p = 14'd4403;
            {7'd119,7'd38}:		p = 14'd4522;
            {7'd119,7'd39}:		p = 14'd4641;
            {7'd119,7'd40}:		p = 14'd4760;
            {7'd119,7'd41}:		p = 14'd4879;
            {7'd119,7'd42}:		p = 14'd4998;
            {7'd119,7'd43}:		p = 14'd5117;
            {7'd119,7'd44}:		p = 14'd5236;
            {7'd119,7'd45}:		p = 14'd5355;
            {7'd119,7'd46}:		p = 14'd5474;
            {7'd119,7'd47}:		p = 14'd5593;
            {7'd119,7'd48}:		p = 14'd5712;
            {7'd119,7'd49}:		p = 14'd5831;
            {7'd119,7'd50}:		p = 14'd5950;
            {7'd119,7'd51}:		p = 14'd6069;
            {7'd119,7'd52}:		p = 14'd6188;
            {7'd119,7'd53}:		p = 14'd6307;
            {7'd119,7'd54}:		p = 14'd6426;
            {7'd119,7'd55}:		p = 14'd6545;
            {7'd119,7'd56}:		p = 14'd6664;
            {7'd119,7'd57}:		p = 14'd6783;
            {7'd119,7'd58}:		p = 14'd6902;
            {7'd119,7'd59}:		p = 14'd7021;
            {7'd119,7'd60}:		p = 14'd7140;
            {7'd119,7'd61}:		p = 14'd7259;
            {7'd119,7'd62}:		p = 14'd7378;
            {7'd119,7'd63}:		p = 14'd7497;
            {7'd119,7'd64}:		p = 14'd7616;
            {7'd119,7'd65}:		p = 14'd7735;
            {7'd119,7'd66}:		p = 14'd7854;
            {7'd119,7'd67}:		p = 14'd7973;
            {7'd119,7'd68}:		p = 14'd8092;
            {7'd119,7'd69}:		p = 14'd8211;
            {7'd119,7'd70}:		p = 14'd8330;
            {7'd119,7'd71}:		p = 14'd8449;
            {7'd119,7'd72}:		p = 14'd8568;
            {7'd119,7'd73}:		p = 14'd8687;
            {7'd119,7'd74}:		p = 14'd8806;
            {7'd119,7'd75}:		p = 14'd8925;
            {7'd119,7'd76}:		p = 14'd9044;
            {7'd119,7'd77}:		p = 14'd9163;
            {7'd119,7'd78}:		p = 14'd9282;
            {7'd119,7'd79}:		p = 14'd9401;
            {7'd119,7'd80}:		p = 14'd9520;
            {7'd119,7'd81}:		p = 14'd9639;
            {7'd119,7'd82}:		p = 14'd9758;
            {7'd119,7'd83}:		p = 14'd9877;
            {7'd119,7'd84}:		p = 14'd9996;
            {7'd119,7'd85}:		p = 14'd10115;
            {7'd119,7'd86}:		p = 14'd10234;
            {7'd119,7'd87}:		p = 14'd10353;
            {7'd119,7'd88}:		p = 14'd10472;
            {7'd119,7'd89}:		p = 14'd10591;
            {7'd119,7'd90}:		p = 14'd10710;
            {7'd119,7'd91}:		p = 14'd10829;
            {7'd119,7'd92}:		p = 14'd10948;
            {7'd119,7'd93}:		p = 14'd11067;
            {7'd119,7'd94}:		p = 14'd11186;
            {7'd119,7'd95}:		p = 14'd11305;
            {7'd119,7'd96}:		p = 14'd11424;
            {7'd119,7'd97}:		p = 14'd11543;
            {7'd119,7'd98}:		p = 14'd11662;
            {7'd119,7'd99}:		p = 14'd11781;
            {7'd119,7'd100}:		p = 14'd11900;
            {7'd119,7'd101}:		p = 14'd12019;
            {7'd119,7'd102}:		p = 14'd12138;
            {7'd119,7'd103}:		p = 14'd12257;
            {7'd119,7'd104}:		p = 14'd12376;
            {7'd119,7'd105}:		p = 14'd12495;
            {7'd119,7'd106}:		p = 14'd12614;
            {7'd119,7'd107}:		p = 14'd12733;
            {7'd119,7'd108}:		p = 14'd12852;
            {7'd119,7'd109}:		p = 14'd12971;
            {7'd119,7'd110}:		p = 14'd13090;
            {7'd119,7'd111}:		p = 14'd13209;
            {7'd119,7'd112}:		p = 14'd13328;
            {7'd119,7'd113}:		p = 14'd13447;
            {7'd119,7'd114}:		p = 14'd13566;
            {7'd119,7'd115}:		p = 14'd13685;
            {7'd119,7'd116}:		p = 14'd13804;
            {7'd119,7'd117}:		p = 14'd13923;
            {7'd119,7'd118}:		p = 14'd14042;
            {7'd119,7'd119}:		p = 14'd14161;
            {7'd119,7'd120}:		p = 14'd14280;
            {7'd119,7'd121}:		p = 14'd14399;
            {7'd119,7'd122}:		p = 14'd14518;
            {7'd119,7'd123}:		p = 14'd14637;
            {7'd119,7'd124}:		p = 14'd14756;
            {7'd119,7'd125}:		p = 14'd14875;
            {7'd119,7'd126}:		p = 14'd14994;
            {7'd119,7'd127}:		p = 14'd15113;
            {7'd120,7'd0}:		p = 14'd0;
            {7'd120,7'd1}:		p = 14'd120;
            {7'd120,7'd2}:		p = 14'd240;
            {7'd120,7'd3}:		p = 14'd360;
            {7'd120,7'd4}:		p = 14'd480;
            {7'd120,7'd5}:		p = 14'd600;
            {7'd120,7'd6}:		p = 14'd720;
            {7'd120,7'd7}:		p = 14'd840;
            {7'd120,7'd8}:		p = 14'd960;
            {7'd120,7'd9}:		p = 14'd1080;
            {7'd120,7'd10}:		p = 14'd1200;
            {7'd120,7'd11}:		p = 14'd1320;
            {7'd120,7'd12}:		p = 14'd1440;
            {7'd120,7'd13}:		p = 14'd1560;
            {7'd120,7'd14}:		p = 14'd1680;
            {7'd120,7'd15}:		p = 14'd1800;
            {7'd120,7'd16}:		p = 14'd1920;
            {7'd120,7'd17}:		p = 14'd2040;
            {7'd120,7'd18}:		p = 14'd2160;
            {7'd120,7'd19}:		p = 14'd2280;
            {7'd120,7'd20}:		p = 14'd2400;
            {7'd120,7'd21}:		p = 14'd2520;
            {7'd120,7'd22}:		p = 14'd2640;
            {7'd120,7'd23}:		p = 14'd2760;
            {7'd120,7'd24}:		p = 14'd2880;
            {7'd120,7'd25}:		p = 14'd3000;
            {7'd120,7'd26}:		p = 14'd3120;
            {7'd120,7'd27}:		p = 14'd3240;
            {7'd120,7'd28}:		p = 14'd3360;
            {7'd120,7'd29}:		p = 14'd3480;
            {7'd120,7'd30}:		p = 14'd3600;
            {7'd120,7'd31}:		p = 14'd3720;
            {7'd120,7'd32}:		p = 14'd3840;
            {7'd120,7'd33}:		p = 14'd3960;
            {7'd120,7'd34}:		p = 14'd4080;
            {7'd120,7'd35}:		p = 14'd4200;
            {7'd120,7'd36}:		p = 14'd4320;
            {7'd120,7'd37}:		p = 14'd4440;
            {7'd120,7'd38}:		p = 14'd4560;
            {7'd120,7'd39}:		p = 14'd4680;
            {7'd120,7'd40}:		p = 14'd4800;
            {7'd120,7'd41}:		p = 14'd4920;
            {7'd120,7'd42}:		p = 14'd5040;
            {7'd120,7'd43}:		p = 14'd5160;
            {7'd120,7'd44}:		p = 14'd5280;
            {7'd120,7'd45}:		p = 14'd5400;
            {7'd120,7'd46}:		p = 14'd5520;
            {7'd120,7'd47}:		p = 14'd5640;
            {7'd120,7'd48}:		p = 14'd5760;
            {7'd120,7'd49}:		p = 14'd5880;
            {7'd120,7'd50}:		p = 14'd6000;
            {7'd120,7'd51}:		p = 14'd6120;
            {7'd120,7'd52}:		p = 14'd6240;
            {7'd120,7'd53}:		p = 14'd6360;
            {7'd120,7'd54}:		p = 14'd6480;
            {7'd120,7'd55}:		p = 14'd6600;
            {7'd120,7'd56}:		p = 14'd6720;
            {7'd120,7'd57}:		p = 14'd6840;
            {7'd120,7'd58}:		p = 14'd6960;
            {7'd120,7'd59}:		p = 14'd7080;
            {7'd120,7'd60}:		p = 14'd7200;
            {7'd120,7'd61}:		p = 14'd7320;
            {7'd120,7'd62}:		p = 14'd7440;
            {7'd120,7'd63}:		p = 14'd7560;
            {7'd120,7'd64}:		p = 14'd7680;
            {7'd120,7'd65}:		p = 14'd7800;
            {7'd120,7'd66}:		p = 14'd7920;
            {7'd120,7'd67}:		p = 14'd8040;
            {7'd120,7'd68}:		p = 14'd8160;
            {7'd120,7'd69}:		p = 14'd8280;
            {7'd120,7'd70}:		p = 14'd8400;
            {7'd120,7'd71}:		p = 14'd8520;
            {7'd120,7'd72}:		p = 14'd8640;
            {7'd120,7'd73}:		p = 14'd8760;
            {7'd120,7'd74}:		p = 14'd8880;
            {7'd120,7'd75}:		p = 14'd9000;
            {7'd120,7'd76}:		p = 14'd9120;
            {7'd120,7'd77}:		p = 14'd9240;
            {7'd120,7'd78}:		p = 14'd9360;
            {7'd120,7'd79}:		p = 14'd9480;
            {7'd120,7'd80}:		p = 14'd9600;
            {7'd120,7'd81}:		p = 14'd9720;
            {7'd120,7'd82}:		p = 14'd9840;
            {7'd120,7'd83}:		p = 14'd9960;
            {7'd120,7'd84}:		p = 14'd10080;
            {7'd120,7'd85}:		p = 14'd10200;
            {7'd120,7'd86}:		p = 14'd10320;
            {7'd120,7'd87}:		p = 14'd10440;
            {7'd120,7'd88}:		p = 14'd10560;
            {7'd120,7'd89}:		p = 14'd10680;
            {7'd120,7'd90}:		p = 14'd10800;
            {7'd120,7'd91}:		p = 14'd10920;
            {7'd120,7'd92}:		p = 14'd11040;
            {7'd120,7'd93}:		p = 14'd11160;
            {7'd120,7'd94}:		p = 14'd11280;
            {7'd120,7'd95}:		p = 14'd11400;
            {7'd120,7'd96}:		p = 14'd11520;
            {7'd120,7'd97}:		p = 14'd11640;
            {7'd120,7'd98}:		p = 14'd11760;
            {7'd120,7'd99}:		p = 14'd11880;
            {7'd120,7'd100}:		p = 14'd12000;
            {7'd120,7'd101}:		p = 14'd12120;
            {7'd120,7'd102}:		p = 14'd12240;
            {7'd120,7'd103}:		p = 14'd12360;
            {7'd120,7'd104}:		p = 14'd12480;
            {7'd120,7'd105}:		p = 14'd12600;
            {7'd120,7'd106}:		p = 14'd12720;
            {7'd120,7'd107}:		p = 14'd12840;
            {7'd120,7'd108}:		p = 14'd12960;
            {7'd120,7'd109}:		p = 14'd13080;
            {7'd120,7'd110}:		p = 14'd13200;
            {7'd120,7'd111}:		p = 14'd13320;
            {7'd120,7'd112}:		p = 14'd13440;
            {7'd120,7'd113}:		p = 14'd13560;
            {7'd120,7'd114}:		p = 14'd13680;
            {7'd120,7'd115}:		p = 14'd13800;
            {7'd120,7'd116}:		p = 14'd13920;
            {7'd120,7'd117}:		p = 14'd14040;
            {7'd120,7'd118}:		p = 14'd14160;
            {7'd120,7'd119}:		p = 14'd14280;
            {7'd120,7'd120}:		p = 14'd14400;
            {7'd120,7'd121}:		p = 14'd14520;
            {7'd120,7'd122}:		p = 14'd14640;
            {7'd120,7'd123}:		p = 14'd14760;
            {7'd120,7'd124}:		p = 14'd14880;
            {7'd120,7'd125}:		p = 14'd15000;
            {7'd120,7'd126}:		p = 14'd15120;
            {7'd120,7'd127}:		p = 14'd15240;
            {7'd121,7'd0}:		p = 14'd0;
            {7'd121,7'd1}:		p = 14'd121;
            {7'd121,7'd2}:		p = 14'd242;
            {7'd121,7'd3}:		p = 14'd363;
            {7'd121,7'd4}:		p = 14'd484;
            {7'd121,7'd5}:		p = 14'd605;
            {7'd121,7'd6}:		p = 14'd726;
            {7'd121,7'd7}:		p = 14'd847;
            {7'd121,7'd8}:		p = 14'd968;
            {7'd121,7'd9}:		p = 14'd1089;
            {7'd121,7'd10}:		p = 14'd1210;
            {7'd121,7'd11}:		p = 14'd1331;
            {7'd121,7'd12}:		p = 14'd1452;
            {7'd121,7'd13}:		p = 14'd1573;
            {7'd121,7'd14}:		p = 14'd1694;
            {7'd121,7'd15}:		p = 14'd1815;
            {7'd121,7'd16}:		p = 14'd1936;
            {7'd121,7'd17}:		p = 14'd2057;
            {7'd121,7'd18}:		p = 14'd2178;
            {7'd121,7'd19}:		p = 14'd2299;
            {7'd121,7'd20}:		p = 14'd2420;
            {7'd121,7'd21}:		p = 14'd2541;
            {7'd121,7'd22}:		p = 14'd2662;
            {7'd121,7'd23}:		p = 14'd2783;
            {7'd121,7'd24}:		p = 14'd2904;
            {7'd121,7'd25}:		p = 14'd3025;
            {7'd121,7'd26}:		p = 14'd3146;
            {7'd121,7'd27}:		p = 14'd3267;
            {7'd121,7'd28}:		p = 14'd3388;
            {7'd121,7'd29}:		p = 14'd3509;
            {7'd121,7'd30}:		p = 14'd3630;
            {7'd121,7'd31}:		p = 14'd3751;
            {7'd121,7'd32}:		p = 14'd3872;
            {7'd121,7'd33}:		p = 14'd3993;
            {7'd121,7'd34}:		p = 14'd4114;
            {7'd121,7'd35}:		p = 14'd4235;
            {7'd121,7'd36}:		p = 14'd4356;
            {7'd121,7'd37}:		p = 14'd4477;
            {7'd121,7'd38}:		p = 14'd4598;
            {7'd121,7'd39}:		p = 14'd4719;
            {7'd121,7'd40}:		p = 14'd4840;
            {7'd121,7'd41}:		p = 14'd4961;
            {7'd121,7'd42}:		p = 14'd5082;
            {7'd121,7'd43}:		p = 14'd5203;
            {7'd121,7'd44}:		p = 14'd5324;
            {7'd121,7'd45}:		p = 14'd5445;
            {7'd121,7'd46}:		p = 14'd5566;
            {7'd121,7'd47}:		p = 14'd5687;
            {7'd121,7'd48}:		p = 14'd5808;
            {7'd121,7'd49}:		p = 14'd5929;
            {7'd121,7'd50}:		p = 14'd6050;
            {7'd121,7'd51}:		p = 14'd6171;
            {7'd121,7'd52}:		p = 14'd6292;
            {7'd121,7'd53}:		p = 14'd6413;
            {7'd121,7'd54}:		p = 14'd6534;
            {7'd121,7'd55}:		p = 14'd6655;
            {7'd121,7'd56}:		p = 14'd6776;
            {7'd121,7'd57}:		p = 14'd6897;
            {7'd121,7'd58}:		p = 14'd7018;
            {7'd121,7'd59}:		p = 14'd7139;
            {7'd121,7'd60}:		p = 14'd7260;
            {7'd121,7'd61}:		p = 14'd7381;
            {7'd121,7'd62}:		p = 14'd7502;
            {7'd121,7'd63}:		p = 14'd7623;
            {7'd121,7'd64}:		p = 14'd7744;
            {7'd121,7'd65}:		p = 14'd7865;
            {7'd121,7'd66}:		p = 14'd7986;
            {7'd121,7'd67}:		p = 14'd8107;
            {7'd121,7'd68}:		p = 14'd8228;
            {7'd121,7'd69}:		p = 14'd8349;
            {7'd121,7'd70}:		p = 14'd8470;
            {7'd121,7'd71}:		p = 14'd8591;
            {7'd121,7'd72}:		p = 14'd8712;
            {7'd121,7'd73}:		p = 14'd8833;
            {7'd121,7'd74}:		p = 14'd8954;
            {7'd121,7'd75}:		p = 14'd9075;
            {7'd121,7'd76}:		p = 14'd9196;
            {7'd121,7'd77}:		p = 14'd9317;
            {7'd121,7'd78}:		p = 14'd9438;
            {7'd121,7'd79}:		p = 14'd9559;
            {7'd121,7'd80}:		p = 14'd9680;
            {7'd121,7'd81}:		p = 14'd9801;
            {7'd121,7'd82}:		p = 14'd9922;
            {7'd121,7'd83}:		p = 14'd10043;
            {7'd121,7'd84}:		p = 14'd10164;
            {7'd121,7'd85}:		p = 14'd10285;
            {7'd121,7'd86}:		p = 14'd10406;
            {7'd121,7'd87}:		p = 14'd10527;
            {7'd121,7'd88}:		p = 14'd10648;
            {7'd121,7'd89}:		p = 14'd10769;
            {7'd121,7'd90}:		p = 14'd10890;
            {7'd121,7'd91}:		p = 14'd11011;
            {7'd121,7'd92}:		p = 14'd11132;
            {7'd121,7'd93}:		p = 14'd11253;
            {7'd121,7'd94}:		p = 14'd11374;
            {7'd121,7'd95}:		p = 14'd11495;
            {7'd121,7'd96}:		p = 14'd11616;
            {7'd121,7'd97}:		p = 14'd11737;
            {7'd121,7'd98}:		p = 14'd11858;
            {7'd121,7'd99}:		p = 14'd11979;
            {7'd121,7'd100}:		p = 14'd12100;
            {7'd121,7'd101}:		p = 14'd12221;
            {7'd121,7'd102}:		p = 14'd12342;
            {7'd121,7'd103}:		p = 14'd12463;
            {7'd121,7'd104}:		p = 14'd12584;
            {7'd121,7'd105}:		p = 14'd12705;
            {7'd121,7'd106}:		p = 14'd12826;
            {7'd121,7'd107}:		p = 14'd12947;
            {7'd121,7'd108}:		p = 14'd13068;
            {7'd121,7'd109}:		p = 14'd13189;
            {7'd121,7'd110}:		p = 14'd13310;
            {7'd121,7'd111}:		p = 14'd13431;
            {7'd121,7'd112}:		p = 14'd13552;
            {7'd121,7'd113}:		p = 14'd13673;
            {7'd121,7'd114}:		p = 14'd13794;
            {7'd121,7'd115}:		p = 14'd13915;
            {7'd121,7'd116}:		p = 14'd14036;
            {7'd121,7'd117}:		p = 14'd14157;
            {7'd121,7'd118}:		p = 14'd14278;
            {7'd121,7'd119}:		p = 14'd14399;
            {7'd121,7'd120}:		p = 14'd14520;
            {7'd121,7'd121}:		p = 14'd14641;
            {7'd121,7'd122}:		p = 14'd14762;
            {7'd121,7'd123}:		p = 14'd14883;
            {7'd121,7'd124}:		p = 14'd15004;
            {7'd121,7'd125}:		p = 14'd15125;
            {7'd121,7'd126}:		p = 14'd15246;
            {7'd121,7'd127}:		p = 14'd15367;
            {7'd122,7'd0}:		p = 14'd0;
            {7'd122,7'd1}:		p = 14'd122;
            {7'd122,7'd2}:		p = 14'd244;
            {7'd122,7'd3}:		p = 14'd366;
            {7'd122,7'd4}:		p = 14'd488;
            {7'd122,7'd5}:		p = 14'd610;
            {7'd122,7'd6}:		p = 14'd732;
            {7'd122,7'd7}:		p = 14'd854;
            {7'd122,7'd8}:		p = 14'd976;
            {7'd122,7'd9}:		p = 14'd1098;
            {7'd122,7'd10}:		p = 14'd1220;
            {7'd122,7'd11}:		p = 14'd1342;
            {7'd122,7'd12}:		p = 14'd1464;
            {7'd122,7'd13}:		p = 14'd1586;
            {7'd122,7'd14}:		p = 14'd1708;
            {7'd122,7'd15}:		p = 14'd1830;
            {7'd122,7'd16}:		p = 14'd1952;
            {7'd122,7'd17}:		p = 14'd2074;
            {7'd122,7'd18}:		p = 14'd2196;
            {7'd122,7'd19}:		p = 14'd2318;
            {7'd122,7'd20}:		p = 14'd2440;
            {7'd122,7'd21}:		p = 14'd2562;
            {7'd122,7'd22}:		p = 14'd2684;
            {7'd122,7'd23}:		p = 14'd2806;
            {7'd122,7'd24}:		p = 14'd2928;
            {7'd122,7'd25}:		p = 14'd3050;
            {7'd122,7'd26}:		p = 14'd3172;
            {7'd122,7'd27}:		p = 14'd3294;
            {7'd122,7'd28}:		p = 14'd3416;
            {7'd122,7'd29}:		p = 14'd3538;
            {7'd122,7'd30}:		p = 14'd3660;
            {7'd122,7'd31}:		p = 14'd3782;
            {7'd122,7'd32}:		p = 14'd3904;
            {7'd122,7'd33}:		p = 14'd4026;
            {7'd122,7'd34}:		p = 14'd4148;
            {7'd122,7'd35}:		p = 14'd4270;
            {7'd122,7'd36}:		p = 14'd4392;
            {7'd122,7'd37}:		p = 14'd4514;
            {7'd122,7'd38}:		p = 14'd4636;
            {7'd122,7'd39}:		p = 14'd4758;
            {7'd122,7'd40}:		p = 14'd4880;
            {7'd122,7'd41}:		p = 14'd5002;
            {7'd122,7'd42}:		p = 14'd5124;
            {7'd122,7'd43}:		p = 14'd5246;
            {7'd122,7'd44}:		p = 14'd5368;
            {7'd122,7'd45}:		p = 14'd5490;
            {7'd122,7'd46}:		p = 14'd5612;
            {7'd122,7'd47}:		p = 14'd5734;
            {7'd122,7'd48}:		p = 14'd5856;
            {7'd122,7'd49}:		p = 14'd5978;
            {7'd122,7'd50}:		p = 14'd6100;
            {7'd122,7'd51}:		p = 14'd6222;
            {7'd122,7'd52}:		p = 14'd6344;
            {7'd122,7'd53}:		p = 14'd6466;
            {7'd122,7'd54}:		p = 14'd6588;
            {7'd122,7'd55}:		p = 14'd6710;
            {7'd122,7'd56}:		p = 14'd6832;
            {7'd122,7'd57}:		p = 14'd6954;
            {7'd122,7'd58}:		p = 14'd7076;
            {7'd122,7'd59}:		p = 14'd7198;
            {7'd122,7'd60}:		p = 14'd7320;
            {7'd122,7'd61}:		p = 14'd7442;
            {7'd122,7'd62}:		p = 14'd7564;
            {7'd122,7'd63}:		p = 14'd7686;
            {7'd122,7'd64}:		p = 14'd7808;
            {7'd122,7'd65}:		p = 14'd7930;
            {7'd122,7'd66}:		p = 14'd8052;
            {7'd122,7'd67}:		p = 14'd8174;
            {7'd122,7'd68}:		p = 14'd8296;
            {7'd122,7'd69}:		p = 14'd8418;
            {7'd122,7'd70}:		p = 14'd8540;
            {7'd122,7'd71}:		p = 14'd8662;
            {7'd122,7'd72}:		p = 14'd8784;
            {7'd122,7'd73}:		p = 14'd8906;
            {7'd122,7'd74}:		p = 14'd9028;
            {7'd122,7'd75}:		p = 14'd9150;
            {7'd122,7'd76}:		p = 14'd9272;
            {7'd122,7'd77}:		p = 14'd9394;
            {7'd122,7'd78}:		p = 14'd9516;
            {7'd122,7'd79}:		p = 14'd9638;
            {7'd122,7'd80}:		p = 14'd9760;
            {7'd122,7'd81}:		p = 14'd9882;
            {7'd122,7'd82}:		p = 14'd10004;
            {7'd122,7'd83}:		p = 14'd10126;
            {7'd122,7'd84}:		p = 14'd10248;
            {7'd122,7'd85}:		p = 14'd10370;
            {7'd122,7'd86}:		p = 14'd10492;
            {7'd122,7'd87}:		p = 14'd10614;
            {7'd122,7'd88}:		p = 14'd10736;
            {7'd122,7'd89}:		p = 14'd10858;
            {7'd122,7'd90}:		p = 14'd10980;
            {7'd122,7'd91}:		p = 14'd11102;
            {7'd122,7'd92}:		p = 14'd11224;
            {7'd122,7'd93}:		p = 14'd11346;
            {7'd122,7'd94}:		p = 14'd11468;
            {7'd122,7'd95}:		p = 14'd11590;
            {7'd122,7'd96}:		p = 14'd11712;
            {7'd122,7'd97}:		p = 14'd11834;
            {7'd122,7'd98}:		p = 14'd11956;
            {7'd122,7'd99}:		p = 14'd12078;
            {7'd122,7'd100}:		p = 14'd12200;
            {7'd122,7'd101}:		p = 14'd12322;
            {7'd122,7'd102}:		p = 14'd12444;
            {7'd122,7'd103}:		p = 14'd12566;
            {7'd122,7'd104}:		p = 14'd12688;
            {7'd122,7'd105}:		p = 14'd12810;
            {7'd122,7'd106}:		p = 14'd12932;
            {7'd122,7'd107}:		p = 14'd13054;
            {7'd122,7'd108}:		p = 14'd13176;
            {7'd122,7'd109}:		p = 14'd13298;
            {7'd122,7'd110}:		p = 14'd13420;
            {7'd122,7'd111}:		p = 14'd13542;
            {7'd122,7'd112}:		p = 14'd13664;
            {7'd122,7'd113}:		p = 14'd13786;
            {7'd122,7'd114}:		p = 14'd13908;
            {7'd122,7'd115}:		p = 14'd14030;
            {7'd122,7'd116}:		p = 14'd14152;
            {7'd122,7'd117}:		p = 14'd14274;
            {7'd122,7'd118}:		p = 14'd14396;
            {7'd122,7'd119}:		p = 14'd14518;
            {7'd122,7'd120}:		p = 14'd14640;
            {7'd122,7'd121}:		p = 14'd14762;
            {7'd122,7'd122}:		p = 14'd14884;
            {7'd122,7'd123}:		p = 14'd15006;
            {7'd122,7'd124}:		p = 14'd15128;
            {7'd122,7'd125}:		p = 14'd15250;
            {7'd122,7'd126}:		p = 14'd15372;
            {7'd122,7'd127}:		p = 14'd15494;
            {7'd123,7'd0}:		p = 14'd0;
            {7'd123,7'd1}:		p = 14'd123;
            {7'd123,7'd2}:		p = 14'd246;
            {7'd123,7'd3}:		p = 14'd369;
            {7'd123,7'd4}:		p = 14'd492;
            {7'd123,7'd5}:		p = 14'd615;
            {7'd123,7'd6}:		p = 14'd738;
            {7'd123,7'd7}:		p = 14'd861;
            {7'd123,7'd8}:		p = 14'd984;
            {7'd123,7'd9}:		p = 14'd1107;
            {7'd123,7'd10}:		p = 14'd1230;
            {7'd123,7'd11}:		p = 14'd1353;
            {7'd123,7'd12}:		p = 14'd1476;
            {7'd123,7'd13}:		p = 14'd1599;
            {7'd123,7'd14}:		p = 14'd1722;
            {7'd123,7'd15}:		p = 14'd1845;
            {7'd123,7'd16}:		p = 14'd1968;
            {7'd123,7'd17}:		p = 14'd2091;
            {7'd123,7'd18}:		p = 14'd2214;
            {7'd123,7'd19}:		p = 14'd2337;
            {7'd123,7'd20}:		p = 14'd2460;
            {7'd123,7'd21}:		p = 14'd2583;
            {7'd123,7'd22}:		p = 14'd2706;
            {7'd123,7'd23}:		p = 14'd2829;
            {7'd123,7'd24}:		p = 14'd2952;
            {7'd123,7'd25}:		p = 14'd3075;
            {7'd123,7'd26}:		p = 14'd3198;
            {7'd123,7'd27}:		p = 14'd3321;
            {7'd123,7'd28}:		p = 14'd3444;
            {7'd123,7'd29}:		p = 14'd3567;
            {7'd123,7'd30}:		p = 14'd3690;
            {7'd123,7'd31}:		p = 14'd3813;
            {7'd123,7'd32}:		p = 14'd3936;
            {7'd123,7'd33}:		p = 14'd4059;
            {7'd123,7'd34}:		p = 14'd4182;
            {7'd123,7'd35}:		p = 14'd4305;
            {7'd123,7'd36}:		p = 14'd4428;
            {7'd123,7'd37}:		p = 14'd4551;
            {7'd123,7'd38}:		p = 14'd4674;
            {7'd123,7'd39}:		p = 14'd4797;
            {7'd123,7'd40}:		p = 14'd4920;
            {7'd123,7'd41}:		p = 14'd5043;
            {7'd123,7'd42}:		p = 14'd5166;
            {7'd123,7'd43}:		p = 14'd5289;
            {7'd123,7'd44}:		p = 14'd5412;
            {7'd123,7'd45}:		p = 14'd5535;
            {7'd123,7'd46}:		p = 14'd5658;
            {7'd123,7'd47}:		p = 14'd5781;
            {7'd123,7'd48}:		p = 14'd5904;
            {7'd123,7'd49}:		p = 14'd6027;
            {7'd123,7'd50}:		p = 14'd6150;
            {7'd123,7'd51}:		p = 14'd6273;
            {7'd123,7'd52}:		p = 14'd6396;
            {7'd123,7'd53}:		p = 14'd6519;
            {7'd123,7'd54}:		p = 14'd6642;
            {7'd123,7'd55}:		p = 14'd6765;
            {7'd123,7'd56}:		p = 14'd6888;
            {7'd123,7'd57}:		p = 14'd7011;
            {7'd123,7'd58}:		p = 14'd7134;
            {7'd123,7'd59}:		p = 14'd7257;
            {7'd123,7'd60}:		p = 14'd7380;
            {7'd123,7'd61}:		p = 14'd7503;
            {7'd123,7'd62}:		p = 14'd7626;
            {7'd123,7'd63}:		p = 14'd7749;
            {7'd123,7'd64}:		p = 14'd7872;
            {7'd123,7'd65}:		p = 14'd7995;
            {7'd123,7'd66}:		p = 14'd8118;
            {7'd123,7'd67}:		p = 14'd8241;
            {7'd123,7'd68}:		p = 14'd8364;
            {7'd123,7'd69}:		p = 14'd8487;
            {7'd123,7'd70}:		p = 14'd8610;
            {7'd123,7'd71}:		p = 14'd8733;
            {7'd123,7'd72}:		p = 14'd8856;
            {7'd123,7'd73}:		p = 14'd8979;
            {7'd123,7'd74}:		p = 14'd9102;
            {7'd123,7'd75}:		p = 14'd9225;
            {7'd123,7'd76}:		p = 14'd9348;
            {7'd123,7'd77}:		p = 14'd9471;
            {7'd123,7'd78}:		p = 14'd9594;
            {7'd123,7'd79}:		p = 14'd9717;
            {7'd123,7'd80}:		p = 14'd9840;
            {7'd123,7'd81}:		p = 14'd9963;
            {7'd123,7'd82}:		p = 14'd10086;
            {7'd123,7'd83}:		p = 14'd10209;
            {7'd123,7'd84}:		p = 14'd10332;
            {7'd123,7'd85}:		p = 14'd10455;
            {7'd123,7'd86}:		p = 14'd10578;
            {7'd123,7'd87}:		p = 14'd10701;
            {7'd123,7'd88}:		p = 14'd10824;
            {7'd123,7'd89}:		p = 14'd10947;
            {7'd123,7'd90}:		p = 14'd11070;
            {7'd123,7'd91}:		p = 14'd11193;
            {7'd123,7'd92}:		p = 14'd11316;
            {7'd123,7'd93}:		p = 14'd11439;
            {7'd123,7'd94}:		p = 14'd11562;
            {7'd123,7'd95}:		p = 14'd11685;
            {7'd123,7'd96}:		p = 14'd11808;
            {7'd123,7'd97}:		p = 14'd11931;
            {7'd123,7'd98}:		p = 14'd12054;
            {7'd123,7'd99}:		p = 14'd12177;
            {7'd123,7'd100}:		p = 14'd12300;
            {7'd123,7'd101}:		p = 14'd12423;
            {7'd123,7'd102}:		p = 14'd12546;
            {7'd123,7'd103}:		p = 14'd12669;
            {7'd123,7'd104}:		p = 14'd12792;
            {7'd123,7'd105}:		p = 14'd12915;
            {7'd123,7'd106}:		p = 14'd13038;
            {7'd123,7'd107}:		p = 14'd13161;
            {7'd123,7'd108}:		p = 14'd13284;
            {7'd123,7'd109}:		p = 14'd13407;
            {7'd123,7'd110}:		p = 14'd13530;
            {7'd123,7'd111}:		p = 14'd13653;
            {7'd123,7'd112}:		p = 14'd13776;
            {7'd123,7'd113}:		p = 14'd13899;
            {7'd123,7'd114}:		p = 14'd14022;
            {7'd123,7'd115}:		p = 14'd14145;
            {7'd123,7'd116}:		p = 14'd14268;
            {7'd123,7'd117}:		p = 14'd14391;
            {7'd123,7'd118}:		p = 14'd14514;
            {7'd123,7'd119}:		p = 14'd14637;
            {7'd123,7'd120}:		p = 14'd14760;
            {7'd123,7'd121}:		p = 14'd14883;
            {7'd123,7'd122}:		p = 14'd15006;
            {7'd123,7'd123}:		p = 14'd15129;
            {7'd123,7'd124}:		p = 14'd15252;
            {7'd123,7'd125}:		p = 14'd15375;
            {7'd123,7'd126}:		p = 14'd15498;
            {7'd123,7'd127}:		p = 14'd15621;
            {7'd124,7'd0}:		p = 14'd0;
            {7'd124,7'd1}:		p = 14'd124;
            {7'd124,7'd2}:		p = 14'd248;
            {7'd124,7'd3}:		p = 14'd372;
            {7'd124,7'd4}:		p = 14'd496;
            {7'd124,7'd5}:		p = 14'd620;
            {7'd124,7'd6}:		p = 14'd744;
            {7'd124,7'd7}:		p = 14'd868;
            {7'd124,7'd8}:		p = 14'd992;
            {7'd124,7'd9}:		p = 14'd1116;
            {7'd124,7'd10}:		p = 14'd1240;
            {7'd124,7'd11}:		p = 14'd1364;
            {7'd124,7'd12}:		p = 14'd1488;
            {7'd124,7'd13}:		p = 14'd1612;
            {7'd124,7'd14}:		p = 14'd1736;
            {7'd124,7'd15}:		p = 14'd1860;
            {7'd124,7'd16}:		p = 14'd1984;
            {7'd124,7'd17}:		p = 14'd2108;
            {7'd124,7'd18}:		p = 14'd2232;
            {7'd124,7'd19}:		p = 14'd2356;
            {7'd124,7'd20}:		p = 14'd2480;
            {7'd124,7'd21}:		p = 14'd2604;
            {7'd124,7'd22}:		p = 14'd2728;
            {7'd124,7'd23}:		p = 14'd2852;
            {7'd124,7'd24}:		p = 14'd2976;
            {7'd124,7'd25}:		p = 14'd3100;
            {7'd124,7'd26}:		p = 14'd3224;
            {7'd124,7'd27}:		p = 14'd3348;
            {7'd124,7'd28}:		p = 14'd3472;
            {7'd124,7'd29}:		p = 14'd3596;
            {7'd124,7'd30}:		p = 14'd3720;
            {7'd124,7'd31}:		p = 14'd3844;
            {7'd124,7'd32}:		p = 14'd3968;
            {7'd124,7'd33}:		p = 14'd4092;
            {7'd124,7'd34}:		p = 14'd4216;
            {7'd124,7'd35}:		p = 14'd4340;
            {7'd124,7'd36}:		p = 14'd4464;
            {7'd124,7'd37}:		p = 14'd4588;
            {7'd124,7'd38}:		p = 14'd4712;
            {7'd124,7'd39}:		p = 14'd4836;
            {7'd124,7'd40}:		p = 14'd4960;
            {7'd124,7'd41}:		p = 14'd5084;
            {7'd124,7'd42}:		p = 14'd5208;
            {7'd124,7'd43}:		p = 14'd5332;
            {7'd124,7'd44}:		p = 14'd5456;
            {7'd124,7'd45}:		p = 14'd5580;
            {7'd124,7'd46}:		p = 14'd5704;
            {7'd124,7'd47}:		p = 14'd5828;
            {7'd124,7'd48}:		p = 14'd5952;
            {7'd124,7'd49}:		p = 14'd6076;
            {7'd124,7'd50}:		p = 14'd6200;
            {7'd124,7'd51}:		p = 14'd6324;
            {7'd124,7'd52}:		p = 14'd6448;
            {7'd124,7'd53}:		p = 14'd6572;
            {7'd124,7'd54}:		p = 14'd6696;
            {7'd124,7'd55}:		p = 14'd6820;
            {7'd124,7'd56}:		p = 14'd6944;
            {7'd124,7'd57}:		p = 14'd7068;
            {7'd124,7'd58}:		p = 14'd7192;
            {7'd124,7'd59}:		p = 14'd7316;
            {7'd124,7'd60}:		p = 14'd7440;
            {7'd124,7'd61}:		p = 14'd7564;
            {7'd124,7'd62}:		p = 14'd7688;
            {7'd124,7'd63}:		p = 14'd7812;
            {7'd124,7'd64}:		p = 14'd7936;
            {7'd124,7'd65}:		p = 14'd8060;
            {7'd124,7'd66}:		p = 14'd8184;
            {7'd124,7'd67}:		p = 14'd8308;
            {7'd124,7'd68}:		p = 14'd8432;
            {7'd124,7'd69}:		p = 14'd8556;
            {7'd124,7'd70}:		p = 14'd8680;
            {7'd124,7'd71}:		p = 14'd8804;
            {7'd124,7'd72}:		p = 14'd8928;
            {7'd124,7'd73}:		p = 14'd9052;
            {7'd124,7'd74}:		p = 14'd9176;
            {7'd124,7'd75}:		p = 14'd9300;
            {7'd124,7'd76}:		p = 14'd9424;
            {7'd124,7'd77}:		p = 14'd9548;
            {7'd124,7'd78}:		p = 14'd9672;
            {7'd124,7'd79}:		p = 14'd9796;
            {7'd124,7'd80}:		p = 14'd9920;
            {7'd124,7'd81}:		p = 14'd10044;
            {7'd124,7'd82}:		p = 14'd10168;
            {7'd124,7'd83}:		p = 14'd10292;
            {7'd124,7'd84}:		p = 14'd10416;
            {7'd124,7'd85}:		p = 14'd10540;
            {7'd124,7'd86}:		p = 14'd10664;
            {7'd124,7'd87}:		p = 14'd10788;
            {7'd124,7'd88}:		p = 14'd10912;
            {7'd124,7'd89}:		p = 14'd11036;
            {7'd124,7'd90}:		p = 14'd11160;
            {7'd124,7'd91}:		p = 14'd11284;
            {7'd124,7'd92}:		p = 14'd11408;
            {7'd124,7'd93}:		p = 14'd11532;
            {7'd124,7'd94}:		p = 14'd11656;
            {7'd124,7'd95}:		p = 14'd11780;
            {7'd124,7'd96}:		p = 14'd11904;
            {7'd124,7'd97}:		p = 14'd12028;
            {7'd124,7'd98}:		p = 14'd12152;
            {7'd124,7'd99}:		p = 14'd12276;
            {7'd124,7'd100}:		p = 14'd12400;
            {7'd124,7'd101}:		p = 14'd12524;
            {7'd124,7'd102}:		p = 14'd12648;
            {7'd124,7'd103}:		p = 14'd12772;
            {7'd124,7'd104}:		p = 14'd12896;
            {7'd124,7'd105}:		p = 14'd13020;
            {7'd124,7'd106}:		p = 14'd13144;
            {7'd124,7'd107}:		p = 14'd13268;
            {7'd124,7'd108}:		p = 14'd13392;
            {7'd124,7'd109}:		p = 14'd13516;
            {7'd124,7'd110}:		p = 14'd13640;
            {7'd124,7'd111}:		p = 14'd13764;
            {7'd124,7'd112}:		p = 14'd13888;
            {7'd124,7'd113}:		p = 14'd14012;
            {7'd124,7'd114}:		p = 14'd14136;
            {7'd124,7'd115}:		p = 14'd14260;
            {7'd124,7'd116}:		p = 14'd14384;
            {7'd124,7'd117}:		p = 14'd14508;
            {7'd124,7'd118}:		p = 14'd14632;
            {7'd124,7'd119}:		p = 14'd14756;
            {7'd124,7'd120}:		p = 14'd14880;
            {7'd124,7'd121}:		p = 14'd15004;
            {7'd124,7'd122}:		p = 14'd15128;
            {7'd124,7'd123}:		p = 14'd15252;
            {7'd124,7'd124}:		p = 14'd15376;
            {7'd124,7'd125}:		p = 14'd15500;
            {7'd124,7'd126}:		p = 14'd15624;
            {7'd124,7'd127}:		p = 14'd15748;
            {7'd125,7'd0}:		p = 14'd0;
            {7'd125,7'd1}:		p = 14'd125;
            {7'd125,7'd2}:		p = 14'd250;
            {7'd125,7'd3}:		p = 14'd375;
            {7'd125,7'd4}:		p = 14'd500;
            {7'd125,7'd5}:		p = 14'd625;
            {7'd125,7'd6}:		p = 14'd750;
            {7'd125,7'd7}:		p = 14'd875;
            {7'd125,7'd8}:		p = 14'd1000;
            {7'd125,7'd9}:		p = 14'd1125;
            {7'd125,7'd10}:		p = 14'd1250;
            {7'd125,7'd11}:		p = 14'd1375;
            {7'd125,7'd12}:		p = 14'd1500;
            {7'd125,7'd13}:		p = 14'd1625;
            {7'd125,7'd14}:		p = 14'd1750;
            {7'd125,7'd15}:		p = 14'd1875;
            {7'd125,7'd16}:		p = 14'd2000;
            {7'd125,7'd17}:		p = 14'd2125;
            {7'd125,7'd18}:		p = 14'd2250;
            {7'd125,7'd19}:		p = 14'd2375;
            {7'd125,7'd20}:		p = 14'd2500;
            {7'd125,7'd21}:		p = 14'd2625;
            {7'd125,7'd22}:		p = 14'd2750;
            {7'd125,7'd23}:		p = 14'd2875;
            {7'd125,7'd24}:		p = 14'd3000;
            {7'd125,7'd25}:		p = 14'd3125;
            {7'd125,7'd26}:		p = 14'd3250;
            {7'd125,7'd27}:		p = 14'd3375;
            {7'd125,7'd28}:		p = 14'd3500;
            {7'd125,7'd29}:		p = 14'd3625;
            {7'd125,7'd30}:		p = 14'd3750;
            {7'd125,7'd31}:		p = 14'd3875;
            {7'd125,7'd32}:		p = 14'd4000;
            {7'd125,7'd33}:		p = 14'd4125;
            {7'd125,7'd34}:		p = 14'd4250;
            {7'd125,7'd35}:		p = 14'd4375;
            {7'd125,7'd36}:		p = 14'd4500;
            {7'd125,7'd37}:		p = 14'd4625;
            {7'd125,7'd38}:		p = 14'd4750;
            {7'd125,7'd39}:		p = 14'd4875;
            {7'd125,7'd40}:		p = 14'd5000;
            {7'd125,7'd41}:		p = 14'd5125;
            {7'd125,7'd42}:		p = 14'd5250;
            {7'd125,7'd43}:		p = 14'd5375;
            {7'd125,7'd44}:		p = 14'd5500;
            {7'd125,7'd45}:		p = 14'd5625;
            {7'd125,7'd46}:		p = 14'd5750;
            {7'd125,7'd47}:		p = 14'd5875;
            {7'd125,7'd48}:		p = 14'd6000;
            {7'd125,7'd49}:		p = 14'd6125;
            {7'd125,7'd50}:		p = 14'd6250;
            {7'd125,7'd51}:		p = 14'd6375;
            {7'd125,7'd52}:		p = 14'd6500;
            {7'd125,7'd53}:		p = 14'd6625;
            {7'd125,7'd54}:		p = 14'd6750;
            {7'd125,7'd55}:		p = 14'd6875;
            {7'd125,7'd56}:		p = 14'd7000;
            {7'd125,7'd57}:		p = 14'd7125;
            {7'd125,7'd58}:		p = 14'd7250;
            {7'd125,7'd59}:		p = 14'd7375;
            {7'd125,7'd60}:		p = 14'd7500;
            {7'd125,7'd61}:		p = 14'd7625;
            {7'd125,7'd62}:		p = 14'd7750;
            {7'd125,7'd63}:		p = 14'd7875;
            {7'd125,7'd64}:		p = 14'd8000;
            {7'd125,7'd65}:		p = 14'd8125;
            {7'd125,7'd66}:		p = 14'd8250;
            {7'd125,7'd67}:		p = 14'd8375;
            {7'd125,7'd68}:		p = 14'd8500;
            {7'd125,7'd69}:		p = 14'd8625;
            {7'd125,7'd70}:		p = 14'd8750;
            {7'd125,7'd71}:		p = 14'd8875;
            {7'd125,7'd72}:		p = 14'd9000;
            {7'd125,7'd73}:		p = 14'd9125;
            {7'd125,7'd74}:		p = 14'd9250;
            {7'd125,7'd75}:		p = 14'd9375;
            {7'd125,7'd76}:		p = 14'd9500;
            {7'd125,7'd77}:		p = 14'd9625;
            {7'd125,7'd78}:		p = 14'd9750;
            {7'd125,7'd79}:		p = 14'd9875;
            {7'd125,7'd80}:		p = 14'd10000;
            {7'd125,7'd81}:		p = 14'd10125;
            {7'd125,7'd82}:		p = 14'd10250;
            {7'd125,7'd83}:		p = 14'd10375;
            {7'd125,7'd84}:		p = 14'd10500;
            {7'd125,7'd85}:		p = 14'd10625;
            {7'd125,7'd86}:		p = 14'd10750;
            {7'd125,7'd87}:		p = 14'd10875;
            {7'd125,7'd88}:		p = 14'd11000;
            {7'd125,7'd89}:		p = 14'd11125;
            {7'd125,7'd90}:		p = 14'd11250;
            {7'd125,7'd91}:		p = 14'd11375;
            {7'd125,7'd92}:		p = 14'd11500;
            {7'd125,7'd93}:		p = 14'd11625;
            {7'd125,7'd94}:		p = 14'd11750;
            {7'd125,7'd95}:		p = 14'd11875;
            {7'd125,7'd96}:		p = 14'd12000;
            {7'd125,7'd97}:		p = 14'd12125;
            {7'd125,7'd98}:		p = 14'd12250;
            {7'd125,7'd99}:		p = 14'd12375;
            {7'd125,7'd100}:		p = 14'd12500;
            {7'd125,7'd101}:		p = 14'd12625;
            {7'd125,7'd102}:		p = 14'd12750;
            {7'd125,7'd103}:		p = 14'd12875;
            {7'd125,7'd104}:		p = 14'd13000;
            {7'd125,7'd105}:		p = 14'd13125;
            {7'd125,7'd106}:		p = 14'd13250;
            {7'd125,7'd107}:		p = 14'd13375;
            {7'd125,7'd108}:		p = 14'd13500;
            {7'd125,7'd109}:		p = 14'd13625;
            {7'd125,7'd110}:		p = 14'd13750;
            {7'd125,7'd111}:		p = 14'd13875;
            {7'd125,7'd112}:		p = 14'd14000;
            {7'd125,7'd113}:		p = 14'd14125;
            {7'd125,7'd114}:		p = 14'd14250;
            {7'd125,7'd115}:		p = 14'd14375;
            {7'd125,7'd116}:		p = 14'd14500;
            {7'd125,7'd117}:		p = 14'd14625;
            {7'd125,7'd118}:		p = 14'd14750;
            {7'd125,7'd119}:		p = 14'd14875;
            {7'd125,7'd120}:		p = 14'd15000;
            {7'd125,7'd121}:		p = 14'd15125;
            {7'd125,7'd122}:		p = 14'd15250;
            {7'd125,7'd123}:		p = 14'd15375;
            {7'd125,7'd124}:		p = 14'd15500;
            {7'd125,7'd125}:		p = 14'd15625;
            {7'd125,7'd126}:		p = 14'd15750;
            {7'd125,7'd127}:		p = 14'd15875;
            {7'd126,7'd0}:		p = 14'd0;
            {7'd126,7'd1}:		p = 14'd126;
            {7'd126,7'd2}:		p = 14'd252;
            {7'd126,7'd3}:		p = 14'd378;
            {7'd126,7'd4}:		p = 14'd504;
            {7'd126,7'd5}:		p = 14'd630;
            {7'd126,7'd6}:		p = 14'd756;
            {7'd126,7'd7}:		p = 14'd882;
            {7'd126,7'd8}:		p = 14'd1008;
            {7'd126,7'd9}:		p = 14'd1134;
            {7'd126,7'd10}:		p = 14'd1260;
            {7'd126,7'd11}:		p = 14'd1386;
            {7'd126,7'd12}:		p = 14'd1512;
            {7'd126,7'd13}:		p = 14'd1638;
            {7'd126,7'd14}:		p = 14'd1764;
            {7'd126,7'd15}:		p = 14'd1890;
            {7'd126,7'd16}:		p = 14'd2016;
            {7'd126,7'd17}:		p = 14'd2142;
            {7'd126,7'd18}:		p = 14'd2268;
            {7'd126,7'd19}:		p = 14'd2394;
            {7'd126,7'd20}:		p = 14'd2520;
            {7'd126,7'd21}:		p = 14'd2646;
            {7'd126,7'd22}:		p = 14'd2772;
            {7'd126,7'd23}:		p = 14'd2898;
            {7'd126,7'd24}:		p = 14'd3024;
            {7'd126,7'd25}:		p = 14'd3150;
            {7'd126,7'd26}:		p = 14'd3276;
            {7'd126,7'd27}:		p = 14'd3402;
            {7'd126,7'd28}:		p = 14'd3528;
            {7'd126,7'd29}:		p = 14'd3654;
            {7'd126,7'd30}:		p = 14'd3780;
            {7'd126,7'd31}:		p = 14'd3906;
            {7'd126,7'd32}:		p = 14'd4032;
            {7'd126,7'd33}:		p = 14'd4158;
            {7'd126,7'd34}:		p = 14'd4284;
            {7'd126,7'd35}:		p = 14'd4410;
            {7'd126,7'd36}:		p = 14'd4536;
            {7'd126,7'd37}:		p = 14'd4662;
            {7'd126,7'd38}:		p = 14'd4788;
            {7'd126,7'd39}:		p = 14'd4914;
            {7'd126,7'd40}:		p = 14'd5040;
            {7'd126,7'd41}:		p = 14'd5166;
            {7'd126,7'd42}:		p = 14'd5292;
            {7'd126,7'd43}:		p = 14'd5418;
            {7'd126,7'd44}:		p = 14'd5544;
            {7'd126,7'd45}:		p = 14'd5670;
            {7'd126,7'd46}:		p = 14'd5796;
            {7'd126,7'd47}:		p = 14'd5922;
            {7'd126,7'd48}:		p = 14'd6048;
            {7'd126,7'd49}:		p = 14'd6174;
            {7'd126,7'd50}:		p = 14'd6300;
            {7'd126,7'd51}:		p = 14'd6426;
            {7'd126,7'd52}:		p = 14'd6552;
            {7'd126,7'd53}:		p = 14'd6678;
            {7'd126,7'd54}:		p = 14'd6804;
            {7'd126,7'd55}:		p = 14'd6930;
            {7'd126,7'd56}:		p = 14'd7056;
            {7'd126,7'd57}:		p = 14'd7182;
            {7'd126,7'd58}:		p = 14'd7308;
            {7'd126,7'd59}:		p = 14'd7434;
            {7'd126,7'd60}:		p = 14'd7560;
            {7'd126,7'd61}:		p = 14'd7686;
            {7'd126,7'd62}:		p = 14'd7812;
            {7'd126,7'd63}:		p = 14'd7938;
            {7'd126,7'd64}:		p = 14'd8064;
            {7'd126,7'd65}:		p = 14'd8190;
            {7'd126,7'd66}:		p = 14'd8316;
            {7'd126,7'd67}:		p = 14'd8442;
            {7'd126,7'd68}:		p = 14'd8568;
            {7'd126,7'd69}:		p = 14'd8694;
            {7'd126,7'd70}:		p = 14'd8820;
            {7'd126,7'd71}:		p = 14'd8946;
            {7'd126,7'd72}:		p = 14'd9072;
            {7'd126,7'd73}:		p = 14'd9198;
            {7'd126,7'd74}:		p = 14'd9324;
            {7'd126,7'd75}:		p = 14'd9450;
            {7'd126,7'd76}:		p = 14'd9576;
            {7'd126,7'd77}:		p = 14'd9702;
            {7'd126,7'd78}:		p = 14'd9828;
            {7'd126,7'd79}:		p = 14'd9954;
            {7'd126,7'd80}:		p = 14'd10080;
            {7'd126,7'd81}:		p = 14'd10206;
            {7'd126,7'd82}:		p = 14'd10332;
            {7'd126,7'd83}:		p = 14'd10458;
            {7'd126,7'd84}:		p = 14'd10584;
            {7'd126,7'd85}:		p = 14'd10710;
            {7'd126,7'd86}:		p = 14'd10836;
            {7'd126,7'd87}:		p = 14'd10962;
            {7'd126,7'd88}:		p = 14'd11088;
            {7'd126,7'd89}:		p = 14'd11214;
            {7'd126,7'd90}:		p = 14'd11340;
            {7'd126,7'd91}:		p = 14'd11466;
            {7'd126,7'd92}:		p = 14'd11592;
            {7'd126,7'd93}:		p = 14'd11718;
            {7'd126,7'd94}:		p = 14'd11844;
            {7'd126,7'd95}:		p = 14'd11970;
            {7'd126,7'd96}:		p = 14'd12096;
            {7'd126,7'd97}:		p = 14'd12222;
            {7'd126,7'd98}:		p = 14'd12348;
            {7'd126,7'd99}:		p = 14'd12474;
            {7'd126,7'd100}:		p = 14'd12600;
            {7'd126,7'd101}:		p = 14'd12726;
            {7'd126,7'd102}:		p = 14'd12852;
            {7'd126,7'd103}:		p = 14'd12978;
            {7'd126,7'd104}:		p = 14'd13104;
            {7'd126,7'd105}:		p = 14'd13230;
            {7'd126,7'd106}:		p = 14'd13356;
            {7'd126,7'd107}:		p = 14'd13482;
            {7'd126,7'd108}:		p = 14'd13608;
            {7'd126,7'd109}:		p = 14'd13734;
            {7'd126,7'd110}:		p = 14'd13860;
            {7'd126,7'd111}:		p = 14'd13986;
            {7'd126,7'd112}:		p = 14'd14112;
            {7'd126,7'd113}:		p = 14'd14238;
            {7'd126,7'd114}:		p = 14'd14364;
            {7'd126,7'd115}:		p = 14'd14490;
            {7'd126,7'd116}:		p = 14'd14616;
            {7'd126,7'd117}:		p = 14'd14742;
            {7'd126,7'd118}:		p = 14'd14868;
            {7'd126,7'd119}:		p = 14'd14994;
            {7'd126,7'd120}:		p = 14'd15120;
            {7'd126,7'd121}:		p = 14'd15246;
            {7'd126,7'd122}:		p = 14'd15372;
            {7'd126,7'd123}:		p = 14'd15498;
            {7'd126,7'd124}:		p = 14'd15624;
            {7'd126,7'd125}:		p = 14'd15750;
            {7'd126,7'd126}:		p = 14'd15876;
            {7'd126,7'd127}:		p = 14'd16002;
            {7'd127,7'd0}:		p = 14'd0;
            {7'd127,7'd1}:		p = 14'd127;
            {7'd127,7'd2}:		p = 14'd254;
            {7'd127,7'd3}:		p = 14'd381;
            {7'd127,7'd4}:		p = 14'd508;
            {7'd127,7'd5}:		p = 14'd635;
            {7'd127,7'd6}:		p = 14'd762;
            {7'd127,7'd7}:		p = 14'd889;
            {7'd127,7'd8}:		p = 14'd1016;
            {7'd127,7'd9}:		p = 14'd1143;
            {7'd127,7'd10}:		p = 14'd1270;
            {7'd127,7'd11}:		p = 14'd1397;
            {7'd127,7'd12}:		p = 14'd1524;
            {7'd127,7'd13}:		p = 14'd1651;
            {7'd127,7'd14}:		p = 14'd1778;
            {7'd127,7'd15}:		p = 14'd1905;
            {7'd127,7'd16}:		p = 14'd2032;
            {7'd127,7'd17}:		p = 14'd2159;
            {7'd127,7'd18}:		p = 14'd2286;
            {7'd127,7'd19}:		p = 14'd2413;
            {7'd127,7'd20}:		p = 14'd2540;
            {7'd127,7'd21}:		p = 14'd2667;
            {7'd127,7'd22}:		p = 14'd2794;
            {7'd127,7'd23}:		p = 14'd2921;
            {7'd127,7'd24}:		p = 14'd3048;
            {7'd127,7'd25}:		p = 14'd3175;
            {7'd127,7'd26}:		p = 14'd3302;
            {7'd127,7'd27}:		p = 14'd3429;
            {7'd127,7'd28}:		p = 14'd3556;
            {7'd127,7'd29}:		p = 14'd3683;
            {7'd127,7'd30}:		p = 14'd3810;
            {7'd127,7'd31}:		p = 14'd3937;
            {7'd127,7'd32}:		p = 14'd4064;
            {7'd127,7'd33}:		p = 14'd4191;
            {7'd127,7'd34}:		p = 14'd4318;
            {7'd127,7'd35}:		p = 14'd4445;
            {7'd127,7'd36}:		p = 14'd4572;
            {7'd127,7'd37}:		p = 14'd4699;
            {7'd127,7'd38}:		p = 14'd4826;
            {7'd127,7'd39}:		p = 14'd4953;
            {7'd127,7'd40}:		p = 14'd5080;
            {7'd127,7'd41}:		p = 14'd5207;
            {7'd127,7'd42}:		p = 14'd5334;
            {7'd127,7'd43}:		p = 14'd5461;
            {7'd127,7'd44}:		p = 14'd5588;
            {7'd127,7'd45}:		p = 14'd5715;
            {7'd127,7'd46}:		p = 14'd5842;
            {7'd127,7'd47}:		p = 14'd5969;
            {7'd127,7'd48}:		p = 14'd6096;
            {7'd127,7'd49}:		p = 14'd6223;
            {7'd127,7'd50}:		p = 14'd6350;
            {7'd127,7'd51}:		p = 14'd6477;
            {7'd127,7'd52}:		p = 14'd6604;
            {7'd127,7'd53}:		p = 14'd6731;
            {7'd127,7'd54}:		p = 14'd6858;
            {7'd127,7'd55}:		p = 14'd6985;
            {7'd127,7'd56}:		p = 14'd7112;
            {7'd127,7'd57}:		p = 14'd7239;
            {7'd127,7'd58}:		p = 14'd7366;
            {7'd127,7'd59}:		p = 14'd7493;
            {7'd127,7'd60}:		p = 14'd7620;
            {7'd127,7'd61}:		p = 14'd7747;
            {7'd127,7'd62}:		p = 14'd7874;
            {7'd127,7'd63}:		p = 14'd8001;
            {7'd127,7'd64}:		p = 14'd8128;
            {7'd127,7'd65}:		p = 14'd8255;
            {7'd127,7'd66}:		p = 14'd8382;
            {7'd127,7'd67}:		p = 14'd8509;
            {7'd127,7'd68}:		p = 14'd8636;
            {7'd127,7'd69}:		p = 14'd8763;
            {7'd127,7'd70}:		p = 14'd8890;
            {7'd127,7'd71}:		p = 14'd9017;
            {7'd127,7'd72}:		p = 14'd9144;
            {7'd127,7'd73}:		p = 14'd9271;
            {7'd127,7'd74}:		p = 14'd9398;
            {7'd127,7'd75}:		p = 14'd9525;
            {7'd127,7'd76}:		p = 14'd9652;
            {7'd127,7'd77}:		p = 14'd9779;
            {7'd127,7'd78}:		p = 14'd9906;
            {7'd127,7'd79}:		p = 14'd10033;
            {7'd127,7'd80}:		p = 14'd10160;
            {7'd127,7'd81}:		p = 14'd10287;
            {7'd127,7'd82}:		p = 14'd10414;
            {7'd127,7'd83}:		p = 14'd10541;
            {7'd127,7'd84}:		p = 14'd10668;
            {7'd127,7'd85}:		p = 14'd10795;
            {7'd127,7'd86}:		p = 14'd10922;
            {7'd127,7'd87}:		p = 14'd11049;
            {7'd127,7'd88}:		p = 14'd11176;
            {7'd127,7'd89}:		p = 14'd11303;
            {7'd127,7'd90}:		p = 14'd11430;
            {7'd127,7'd91}:		p = 14'd11557;
            {7'd127,7'd92}:		p = 14'd11684;
            {7'd127,7'd93}:		p = 14'd11811;
            {7'd127,7'd94}:		p = 14'd11938;
            {7'd127,7'd95}:		p = 14'd12065;
            {7'd127,7'd96}:		p = 14'd12192;
            {7'd127,7'd97}:		p = 14'd12319;
            {7'd127,7'd98}:		p = 14'd12446;
            {7'd127,7'd99}:		p = 14'd12573;
            {7'd127,7'd100}:		p = 14'd12700;
            {7'd127,7'd101}:		p = 14'd12827;
            {7'd127,7'd102}:		p = 14'd12954;
            {7'd127,7'd103}:		p = 14'd13081;
            {7'd127,7'd104}:		p = 14'd13208;
            {7'd127,7'd105}:		p = 14'd13335;
            {7'd127,7'd106}:		p = 14'd13462;
            {7'd127,7'd107}:		p = 14'd13589;
            {7'd127,7'd108}:		p = 14'd13716;
            {7'd127,7'd109}:		p = 14'd13843;
            {7'd127,7'd110}:		p = 14'd13970;
            {7'd127,7'd111}:		p = 14'd14097;
            {7'd127,7'd112}:		p = 14'd14224;
            {7'd127,7'd113}:		p = 14'd14351;
            {7'd127,7'd114}:		p = 14'd14478;
            {7'd127,7'd115}:		p = 14'd14605;
            {7'd127,7'd116}:		p = 14'd14732;
            {7'd127,7'd117}:		p = 14'd14859;
            {7'd127,7'd118}:		p = 14'd14986;
            {7'd127,7'd119}:		p = 14'd15113;
            {7'd127,7'd120}:		p = 14'd15240;
            {7'd127,7'd121}:		p = 14'd15367;
            {7'd127,7'd122}:		p = 14'd15494;
            {7'd127,7'd123}:		p = 14'd15621;
            {7'd127,7'd124}:		p = 14'd15748;
            {7'd127,7'd125}:		p = 14'd15875;
            {7'd127,7'd126}:		p = 14'd16002;
            {7'd127,7'd127}:		p = 14'd16129;
        endcase
    end

//    always_comb begin
//        case (mq)
//            {7'd0,7'd0}:	p <= 14'd0;
//            {7'd0,7'd1}:	p <= 14'd0;
//            14'{7'1,7'1}:	p <= 14'b1;
//            default:       	p <= ~14'd0;
//        endcase
//    end

`ifdef BAR
    //////// FULL ADDERS (RIPPLE CARRY)

    wire [Y_WIDTH-1:0] sum [X_WIDTH-1:0];
    wire [X_WIDTH:0] carry;	// +1

// reg  [(WIDTH<<1)-1:0] add_a[WIDTH-1:0];
// reg  [(WIDTH<<1)-1:0] add_b[WIDTH-1:0];
// wire [(WIDTH<<1)-1:0] add_y[WIDTH-1:0];
//add_a[j] = c;
//add_b[j] = (tmp << j);
//c = add_y[j];	// sum

    assign carry[0] = 0;
    assign sum[0][X_WIDTH-1:0] = { {X_WIDTH-2 {1'b0}}, pp[0][0] };

    genvar piq;
    generate //: genp
        for (piq = 1; piq < Y_WIDTH; piq = piq + 1) begin			// loop 13 times, from 1
            fulladder #(
                .WIDTH(X_WIDTH)
            ) fa (
                .a  (sum[piq-1]),
                .b  (pp[piq] << piq),
                .y  (carry[piq-1]),
                .c  (carry[piq]),
                .s  (sum[piq])
            );
            assign p[piq] = sum[piq][0];
        end
    endgenerate
    
    assign p[0] = sum[0];				// alias for pp[0][0];
    assign p[P_WIDTH-1] = carry[X_WIDTH];		// last carry-out
`endif

`ifdef FOO
    //////// HALF ADDERS

    // adder-sum (alias for final output product)
    //    the LSB (PP0[0]) and MSB (last carry-out) have special treatment
    wire [P_WIDTH-1:0] ads;

    assign ads[0] = pp[0][0];			// LSB output (LSB of PP0 as-is)

    // adder-carry chain
    wire [X_WIDTH:0] acc;			// +1

    // we set this up in preparation for the generate block to cascade
    assign acc[0] = pp[0][1];	// adder-carry maybe this should be external for cascade when supported ?

    // note we start at bit1 as LSB(bit0) has already had special treatment
    generate //: genad
        for(genvar adiq = 1; adiq < Y_WIDTH; adiq++) begin : iq			// loop 1 time, from 1
            for(genvar adim = 1; adim <= X_WIDTH; adim++) begin : im			// loop 2 times, from 1
//                for(genvar adip = adim + 1; adip < adim + 3; adip++) begin : ip	// vanity loop 1 time, from adim + 1
                    // The vanity for loop exists to demonstrate the arcane limitations of verilog :)
                    // In wanting to name my component for better schematic/netlist reading by humans
                    //  adip represents the P (product) output bit we are working on here
                    halfadder #(
                        .WIDTH(1)
                    ) ha (	// ha_$adiq_$adim_$adip => ha_iq1_im1_ip1 ?
                        .a  (acc[adim-1]),
                        .b  (pp[adiq][adim-1]),
                        .s  (ads[adim]),
                        .c  (acc[adim])
                    );
//                end
            end
        end
    endgenerate

    // The generate : genad, above unrolls to look like this:

    // halfadder #(.WIDTH(1)) ha_iq1_im1_ip1
    // (
    //                 .a  (acc[0]),   //(acc[adim-1]),
    //                 .b  (pp[1][0]), //(pp[adiq][adim-1]),
    //                 .s  (ads[1]),   //(ads[adim]),
    //                 .c  (acc[1])    //(acc[adim])
    // );
    // halfadder #(.WIDTH(1)) ha_iq1_im2_ip2
    // (
    //                 .a  (acc[1]),   //(acc[adim-1]),
    //                 .b  (pp[1][1]), //(pp[adiq][adim-1]),
    //                 .s  (ads[2]),   //(acc[adim])
    //                 .c  (acc[2])    //(acc[adim])
    // );

    assign ads[P_WIDTH-1] = acc[X_WIDTH];	// MSB output

    // So this but become easy to see the product
    assign p = ads;
`endif

endmodule
