
`define INPUT_WIDTH	8
`define OUTPUT_WIDTH	8

//`define HAS_SIGN	0
//`define HAS_READY	0

`define READY_FALSE	1'b0
`define READY_TRUE	1'b1
