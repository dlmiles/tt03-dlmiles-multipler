// headline config
`define ONES_WIDTH	4

// wire [7:0] io_in, interface
`define I_CLK_BITID	0
`define I_RST_BITID	1
`define I_I0_BITID	2

// wire [7:0] io_out, interface
`define O_O0_BITID	2
