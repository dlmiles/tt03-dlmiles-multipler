
`define	IMPL_MULU_M7Q7		1
